magic
tech sky130A
magscale 1 2
timestamp 1738263620
<< nwell >>
rect -38 261 1418 582
<< pwell >>
rect 98 157 1318 203
rect 1 21 1318 157
rect 30 -17 64 21
<< locali >>
rect 22 215 88 255
rect 646 323 712 493
rect 814 323 880 493
rect 982 323 1048 493
rect 1150 323 1216 493
rect 646 289 1363 323
rect 1287 181 1363 289
rect 646 147 1363 181
rect 646 52 712 147
rect 814 52 880 147
rect 982 52 1048 147
rect 1150 52 1216 147
<< obsli1 >>
rect 0 527 1380 561
rect 19 323 85 432
rect 119 357 153 527
rect 19 289 156 323
rect 200 309 276 493
rect 122 265 156 289
rect 122 199 208 265
rect 242 255 276 309
rect 310 323 376 493
rect 410 357 444 527
rect 478 323 544 493
rect 578 357 612 527
rect 746 367 780 527
rect 914 367 948 527
rect 1082 367 1116 527
rect 1250 367 1284 527
rect 310 289 612 323
rect 578 255 612 289
rect 242 215 544 255
rect 578 215 1072 255
rect 122 181 156 199
rect 19 147 156 181
rect 242 165 276 215
rect 578 181 612 215
rect 19 52 85 147
rect 119 17 153 113
rect 200 52 276 165
rect 310 147 612 181
rect 310 52 376 147
rect 410 17 444 113
rect 478 52 544 147
rect 578 17 612 113
rect 746 17 780 113
rect 914 17 948 113
rect 1082 17 1116 113
rect 1250 17 1284 113
rect 0 -17 1380 17
<< metal1 >>
rect 0 496 1380 592
rect 0 -48 1380 48
<< labels >>
rlabel locali s 22 215 88 255 6 A
port 1 nsew signal input
rlabel metal1 s 0 -48 1380 48 8 VGND
port 2 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 3 nsew ground bidirectional
rlabel pwell s 1 21 1318 157 6 VNB
port 3 nsew ground bidirectional
rlabel pwell s 98 157 1318 203 6 VNB
port 3 nsew ground bidirectional
rlabel nwell s -38 261 1418 582 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 496 1380 592 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 1150 52 1216 147 6 X
port 6 nsew signal output
rlabel locali s 982 52 1048 147 6 X
port 6 nsew signal output
rlabel locali s 814 52 880 147 6 X
port 6 nsew signal output
rlabel locali s 646 52 712 147 6 X
port 6 nsew signal output
rlabel locali s 646 147 1363 181 6 X
port 6 nsew signal output
rlabel locali s 1287 181 1363 289 6 X
port 6 nsew signal output
rlabel locali s 646 289 1363 323 6 X
port 6 nsew signal output
rlabel locali s 1150 323 1216 493 6 X
port 6 nsew signal output
rlabel locali s 982 323 1048 493 6 X
port 6 nsew signal output
rlabel locali s 814 323 880 493 6 X
port 6 nsew signal output
rlabel locali s 646 323 712 493 6 X
port 6 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1380 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3210828
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3200356
<< end >>
