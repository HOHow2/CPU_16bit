magic
tech sky130A
magscale 1 2
timestamp 1738263620
<< nwell >>
rect -38 261 1510 582
<< pwell >>
rect 1 21 1471 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 415 47 445 177
rect 499 47 529 177
rect 583 47 613 177
rect 667 47 697 177
rect 751 47 781 177
rect 835 47 865 177
rect 919 47 949 177
rect 1003 47 1033 177
rect 1087 47 1117 177
rect 1171 47 1201 177
rect 1255 47 1285 177
rect 1339 47 1369 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 331 297 361 497
rect 415 297 445 497
rect 499 297 529 497
rect 583 297 613 497
rect 667 297 697 497
rect 751 297 781 497
rect 835 297 865 497
rect 919 297 949 497
rect 1003 297 1033 497
rect 1087 297 1117 497
rect 1171 297 1201 497
rect 1255 297 1285 497
rect 1339 297 1369 497
<< ndiff >>
rect 27 165 79 177
rect 27 131 35 165
rect 69 131 79 165
rect 27 97 79 131
rect 27 63 35 97
rect 69 63 79 97
rect 27 47 79 63
rect 109 97 163 177
rect 109 63 119 97
rect 153 63 163 97
rect 109 47 163 63
rect 193 165 247 177
rect 193 131 203 165
rect 237 131 247 165
rect 193 97 247 131
rect 193 63 203 97
rect 237 63 247 97
rect 193 47 247 63
rect 277 97 331 177
rect 277 63 287 97
rect 321 63 331 97
rect 277 47 331 63
rect 361 165 415 177
rect 361 131 371 165
rect 405 131 415 165
rect 361 97 415 131
rect 361 63 371 97
rect 405 63 415 97
rect 361 47 415 63
rect 445 97 499 177
rect 445 63 455 97
rect 489 63 499 97
rect 445 47 499 63
rect 529 165 583 177
rect 529 131 539 165
rect 573 131 583 165
rect 529 97 583 131
rect 529 63 539 97
rect 573 63 583 97
rect 529 47 583 63
rect 613 97 667 177
rect 613 63 623 97
rect 657 63 667 97
rect 613 47 667 63
rect 697 165 751 177
rect 697 131 707 165
rect 741 131 751 165
rect 697 97 751 131
rect 697 63 707 97
rect 741 63 751 97
rect 697 47 751 63
rect 781 165 835 177
rect 781 131 791 165
rect 825 131 835 165
rect 781 47 835 131
rect 865 97 919 177
rect 865 63 875 97
rect 909 63 919 97
rect 865 47 919 63
rect 949 165 1003 177
rect 949 131 959 165
rect 993 131 1003 165
rect 949 47 1003 131
rect 1033 97 1087 177
rect 1033 63 1043 97
rect 1077 63 1087 97
rect 1033 47 1087 63
rect 1117 165 1171 177
rect 1117 131 1127 165
rect 1161 131 1171 165
rect 1117 47 1171 131
rect 1201 97 1255 177
rect 1201 63 1211 97
rect 1245 63 1255 97
rect 1201 47 1255 63
rect 1285 165 1339 177
rect 1285 131 1295 165
rect 1329 131 1339 165
rect 1285 47 1339 131
rect 1369 165 1445 177
rect 1369 131 1399 165
rect 1433 131 1445 165
rect 1369 97 1445 131
rect 1369 63 1399 97
rect 1433 63 1445 97
rect 1369 47 1445 63
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 349 79 383
rect 27 315 35 349
rect 69 315 79 349
rect 27 297 79 315
rect 109 485 163 497
rect 109 451 119 485
rect 153 451 163 485
rect 109 417 163 451
rect 109 383 119 417
rect 153 383 163 417
rect 109 349 163 383
rect 109 315 119 349
rect 153 315 163 349
rect 109 297 163 315
rect 193 485 247 497
rect 193 451 203 485
rect 237 451 247 485
rect 193 417 247 451
rect 193 383 203 417
rect 237 383 247 417
rect 193 297 247 383
rect 277 485 331 497
rect 277 451 287 485
rect 321 451 331 485
rect 277 417 331 451
rect 277 383 287 417
rect 321 383 331 417
rect 277 349 331 383
rect 277 315 287 349
rect 321 315 331 349
rect 277 297 331 315
rect 361 485 415 497
rect 361 451 371 485
rect 405 451 415 485
rect 361 417 415 451
rect 361 383 371 417
rect 405 383 415 417
rect 361 297 415 383
rect 445 485 499 497
rect 445 451 455 485
rect 489 451 499 485
rect 445 417 499 451
rect 445 383 455 417
rect 489 383 499 417
rect 445 349 499 383
rect 445 315 455 349
rect 489 315 499 349
rect 445 297 499 315
rect 529 485 583 497
rect 529 451 539 485
rect 573 451 583 485
rect 529 417 583 451
rect 529 383 539 417
rect 573 383 583 417
rect 529 297 583 383
rect 613 485 667 497
rect 613 451 623 485
rect 657 451 667 485
rect 613 417 667 451
rect 613 383 623 417
rect 657 383 667 417
rect 613 349 667 383
rect 613 315 623 349
rect 657 315 667 349
rect 613 297 667 315
rect 697 485 751 497
rect 697 451 707 485
rect 741 451 751 485
rect 697 417 751 451
rect 697 383 707 417
rect 741 383 751 417
rect 697 297 751 383
rect 781 485 835 497
rect 781 451 791 485
rect 825 451 835 485
rect 781 417 835 451
rect 781 383 791 417
rect 825 383 835 417
rect 781 349 835 383
rect 781 315 791 349
rect 825 315 835 349
rect 781 297 835 315
rect 865 485 919 497
rect 865 451 875 485
rect 909 451 919 485
rect 865 417 919 451
rect 865 383 875 417
rect 909 383 919 417
rect 865 297 919 383
rect 949 485 1003 497
rect 949 451 959 485
rect 993 451 1003 485
rect 949 417 1003 451
rect 949 383 959 417
rect 993 383 1003 417
rect 949 349 1003 383
rect 949 315 959 349
rect 993 315 1003 349
rect 949 297 1003 315
rect 1033 485 1087 497
rect 1033 451 1043 485
rect 1077 451 1087 485
rect 1033 417 1087 451
rect 1033 383 1043 417
rect 1077 383 1087 417
rect 1033 297 1087 383
rect 1117 485 1171 497
rect 1117 451 1127 485
rect 1161 451 1171 485
rect 1117 417 1171 451
rect 1117 383 1127 417
rect 1161 383 1171 417
rect 1117 349 1171 383
rect 1117 315 1127 349
rect 1161 315 1171 349
rect 1117 297 1171 315
rect 1201 485 1255 497
rect 1201 451 1211 485
rect 1245 451 1255 485
rect 1201 417 1255 451
rect 1201 383 1211 417
rect 1245 383 1255 417
rect 1201 297 1255 383
rect 1285 485 1339 497
rect 1285 451 1295 485
rect 1329 451 1339 485
rect 1285 417 1339 451
rect 1285 383 1295 417
rect 1329 383 1339 417
rect 1285 349 1339 383
rect 1285 315 1295 349
rect 1329 315 1339 349
rect 1285 297 1339 315
rect 1369 485 1445 497
rect 1369 451 1399 485
rect 1433 451 1445 485
rect 1369 417 1445 451
rect 1369 383 1399 417
rect 1433 383 1445 417
rect 1369 349 1445 383
rect 1369 315 1399 349
rect 1433 315 1445 349
rect 1369 297 1445 315
<< ndiffc >>
rect 35 131 69 165
rect 35 63 69 97
rect 119 63 153 97
rect 203 131 237 165
rect 203 63 237 97
rect 287 63 321 97
rect 371 131 405 165
rect 371 63 405 97
rect 455 63 489 97
rect 539 131 573 165
rect 539 63 573 97
rect 623 63 657 97
rect 707 131 741 165
rect 707 63 741 97
rect 791 131 825 165
rect 875 63 909 97
rect 959 131 993 165
rect 1043 63 1077 97
rect 1127 131 1161 165
rect 1211 63 1245 97
rect 1295 131 1329 165
rect 1399 131 1433 165
rect 1399 63 1433 97
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 119 451 153 485
rect 119 383 153 417
rect 119 315 153 349
rect 203 451 237 485
rect 203 383 237 417
rect 287 451 321 485
rect 287 383 321 417
rect 287 315 321 349
rect 371 451 405 485
rect 371 383 405 417
rect 455 451 489 485
rect 455 383 489 417
rect 455 315 489 349
rect 539 451 573 485
rect 539 383 573 417
rect 623 451 657 485
rect 623 383 657 417
rect 623 315 657 349
rect 707 451 741 485
rect 707 383 741 417
rect 791 451 825 485
rect 791 383 825 417
rect 791 315 825 349
rect 875 451 909 485
rect 875 383 909 417
rect 959 451 993 485
rect 959 383 993 417
rect 959 315 993 349
rect 1043 451 1077 485
rect 1043 383 1077 417
rect 1127 451 1161 485
rect 1127 383 1161 417
rect 1127 315 1161 349
rect 1211 451 1245 485
rect 1211 383 1245 417
rect 1295 451 1329 485
rect 1295 383 1329 417
rect 1295 315 1329 349
rect 1399 451 1433 485
rect 1399 383 1433 417
rect 1399 315 1433 349
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 331 497 361 523
rect 415 497 445 523
rect 499 497 529 523
rect 583 497 613 523
rect 667 497 697 523
rect 751 497 781 523
rect 835 497 865 523
rect 919 497 949 523
rect 1003 497 1033 523
rect 1087 497 1117 523
rect 1171 497 1201 523
rect 1255 497 1285 523
rect 1339 497 1369 523
rect 79 259 109 297
rect 163 259 193 297
rect 247 259 277 297
rect 331 259 361 297
rect 415 259 445 297
rect 499 259 529 297
rect 583 259 613 297
rect 667 259 697 297
rect 79 249 697 259
rect 79 215 118 249
rect 152 215 203 249
rect 237 215 287 249
rect 321 215 371 249
rect 405 215 455 249
rect 489 215 539 249
rect 573 215 623 249
rect 657 215 697 249
rect 79 205 697 215
rect 79 177 109 205
rect 163 177 193 205
rect 247 177 277 205
rect 331 177 361 205
rect 415 177 445 205
rect 499 177 529 205
rect 583 177 613 205
rect 667 177 697 205
rect 751 259 781 297
rect 835 259 865 297
rect 919 259 949 297
rect 1003 259 1033 297
rect 1087 259 1117 297
rect 1171 259 1201 297
rect 1255 259 1285 297
rect 1339 259 1369 297
rect 751 249 1369 259
rect 751 215 875 249
rect 909 215 959 249
rect 993 215 1043 249
rect 1077 215 1127 249
rect 1161 215 1211 249
rect 1245 215 1369 249
rect 751 205 1369 215
rect 751 177 781 205
rect 835 177 865 205
rect 919 177 949 205
rect 1003 177 1033 205
rect 1087 177 1117 205
rect 1171 177 1201 205
rect 1255 177 1285 205
rect 1339 177 1369 205
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 415 21 445 47
rect 499 21 529 47
rect 583 21 613 47
rect 667 21 697 47
rect 751 21 781 47
rect 835 21 865 47
rect 919 21 949 47
rect 1003 21 1033 47
rect 1087 21 1117 47
rect 1171 21 1201 47
rect 1255 21 1285 47
rect 1339 21 1369 47
<< polycont >>
rect 118 215 152 249
rect 203 215 237 249
rect 287 215 321 249
rect 371 215 405 249
rect 455 215 489 249
rect 539 215 573 249
rect 623 215 657 249
rect 875 215 909 249
rect 959 215 993 249
rect 1043 215 1077 249
rect 1127 215 1161 249
rect 1211 215 1245 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 18 485 69 527
rect 18 451 35 485
rect 18 417 69 451
rect 18 383 35 417
rect 18 349 69 383
rect 18 315 35 349
rect 18 299 69 315
rect 103 485 169 493
rect 103 451 119 485
rect 153 451 169 485
rect 103 417 169 451
rect 103 383 119 417
rect 153 383 169 417
rect 103 349 169 383
rect 203 485 237 527
rect 203 417 237 451
rect 203 367 237 383
rect 271 485 337 493
rect 271 451 287 485
rect 321 451 337 485
rect 271 417 337 451
rect 271 383 287 417
rect 321 383 337 417
rect 103 315 119 349
rect 153 333 169 349
rect 271 349 337 383
rect 371 485 405 527
rect 371 417 405 451
rect 371 367 405 383
rect 439 485 505 493
rect 439 451 455 485
rect 489 451 505 485
rect 439 417 505 451
rect 439 383 455 417
rect 489 383 505 417
rect 271 333 287 349
rect 153 315 287 333
rect 321 333 337 349
rect 439 349 505 383
rect 539 485 573 527
rect 539 417 573 451
rect 539 367 573 383
rect 607 485 673 493
rect 607 451 623 485
rect 657 451 673 485
rect 607 417 673 451
rect 607 383 623 417
rect 657 383 673 417
rect 439 333 455 349
rect 321 315 455 333
rect 489 333 505 349
rect 607 349 673 383
rect 707 485 741 527
rect 707 417 741 451
rect 707 367 741 383
rect 775 485 841 493
rect 775 451 791 485
rect 825 451 841 485
rect 775 417 841 451
rect 775 383 791 417
rect 825 383 841 417
rect 607 333 623 349
rect 489 315 623 333
rect 657 333 673 349
rect 775 349 841 383
rect 875 485 909 527
rect 875 417 909 451
rect 875 367 909 383
rect 943 485 1009 493
rect 943 451 959 485
rect 993 451 1009 485
rect 943 417 1009 451
rect 943 383 959 417
rect 993 383 1009 417
rect 775 333 791 349
rect 657 315 791 333
rect 825 333 841 349
rect 943 349 1009 383
rect 1043 485 1077 527
rect 1043 417 1077 451
rect 1043 367 1077 383
rect 1111 485 1177 493
rect 1111 451 1127 485
rect 1161 451 1177 485
rect 1111 417 1177 451
rect 1111 383 1127 417
rect 1161 383 1177 417
rect 943 333 959 349
rect 825 315 959 333
rect 993 333 1009 349
rect 1111 349 1177 383
rect 1211 485 1245 527
rect 1211 417 1245 451
rect 1211 367 1245 383
rect 1279 485 1345 493
rect 1279 451 1295 485
rect 1329 451 1345 485
rect 1279 417 1345 451
rect 1279 383 1295 417
rect 1329 383 1345 417
rect 1111 333 1127 349
rect 993 315 1127 333
rect 1161 333 1177 349
rect 1279 349 1345 383
rect 1279 333 1295 349
rect 1161 315 1295 333
rect 1329 315 1345 349
rect 103 293 1345 315
rect 1383 485 1454 527
rect 1383 451 1399 485
rect 1433 451 1454 485
rect 1383 417 1454 451
rect 1383 383 1399 417
rect 1433 383 1454 417
rect 1383 349 1454 383
rect 1383 315 1399 349
rect 1433 315 1454 349
rect 1383 299 1454 315
rect 102 249 673 259
rect 102 215 118 249
rect 152 215 203 249
rect 237 215 287 249
rect 321 215 371 249
rect 405 215 455 249
rect 489 215 539 249
rect 573 215 623 249
rect 657 215 673 249
rect 728 215 824 293
rect 858 249 1261 255
rect 858 215 875 249
rect 909 215 959 249
rect 993 215 1043 249
rect 1077 215 1127 249
rect 1161 215 1211 249
rect 1245 215 1261 249
rect 775 181 824 215
rect 1295 181 1345 293
rect 18 165 741 181
rect 18 131 35 165
rect 69 147 203 165
rect 69 131 85 147
rect 18 97 85 131
rect 187 131 203 147
rect 237 147 371 165
rect 237 131 253 147
rect 18 63 35 97
rect 69 63 85 97
rect 18 51 85 63
rect 119 97 153 113
rect 119 17 153 63
rect 187 97 253 131
rect 355 131 371 147
rect 405 147 539 165
rect 405 131 421 147
rect 187 63 203 97
rect 237 63 253 97
rect 187 51 253 63
rect 287 97 321 113
rect 287 17 321 63
rect 355 97 421 131
rect 523 131 539 147
rect 573 147 707 165
rect 573 131 589 147
rect 355 63 371 97
rect 405 63 421 97
rect 355 51 421 63
rect 455 97 489 113
rect 455 17 489 63
rect 523 97 589 131
rect 691 131 707 147
rect 775 165 1345 181
rect 775 131 791 165
rect 825 131 959 165
rect 993 131 1127 165
rect 1161 131 1295 165
rect 1329 131 1345 165
rect 1379 165 1454 181
rect 1379 131 1399 165
rect 1433 131 1454 165
rect 523 63 539 97
rect 573 63 589 97
rect 523 51 589 63
rect 623 97 657 113
rect 623 17 657 63
rect 691 97 741 131
rect 1379 97 1454 131
rect 691 63 707 97
rect 741 63 875 97
rect 909 63 1043 97
rect 1077 63 1211 97
rect 1245 63 1399 97
rect 1433 63 1454 97
rect 691 51 1454 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
<< metal1 >>
rect 0 561 1472 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 0 496 1472 527
rect 0 17 1472 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
rect 0 -48 1472 -17
<< labels >>
flabel locali s 1042 221 1076 255 0 FreeSans 250 0 0 0 A
port 1 nsew signal input
flabel locali s 950 221 984 255 0 FreeSans 250 0 0 0 A
port 1 nsew signal input
flabel locali s 858 221 892 255 0 FreeSans 250 0 0 0 A
port 1 nsew signal input
flabel locali s 582 221 616 255 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel locali s 214 221 248 255 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel locali s 122 221 156 255 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel locali s 766 289 800 323 0 FreeSans 250 0 0 0 Y
port 7 nsew signal output
flabel locali s 766 221 800 255 0 FreeSans 250 0 0 0 Y
port 7 nsew signal output
flabel locali s 1226 221 1260 255 0 FreeSans 250 0 0 0 A
port 1 nsew signal input
flabel locali s 1134 221 1168 255 0 FreeSans 250 0 0 0 A
port 1 nsew signal input
flabel locali s 490 221 524 255 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel locali s 398 221 432 255 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel locali s 306 221 340 255 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 nand2_8
rlabel metal1 s 0 -48 1472 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1472 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1472 544
string GDS_END 1855040
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1842748
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 36.800 0.000 
<< end >>
