magic
tech sky130A
magscale 1 2
timestamp 1738263620
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 532 157 716 203
rect 23 21 716 157
rect 29 -17 63 21
<< locali >>
rect 17 211 155 323
rect 642 299 719 493
rect 663 165 719 299
rect 642 51 719 165
<< obsli1 >>
rect 0 527 736 561
rect 40 401 97 493
rect 131 435 185 527
rect 40 357 231 401
rect 189 177 231 357
rect 40 143 231 177
rect 265 323 345 493
rect 383 401 439 493
rect 543 435 608 527
rect 383 357 608 401
rect 265 211 484 323
rect 518 265 608 357
rect 40 51 97 143
rect 131 17 185 109
rect 265 51 345 211
rect 518 199 629 265
rect 518 177 608 199
rect 383 143 608 177
rect 383 51 439 143
rect 543 17 608 109
rect 0 -17 736 17
<< metal1 >>
rect 0 496 736 592
rect 0 -48 736 48
<< labels >>
rlabel locali s 17 211 155 323 6 A
port 1 nsew signal input
rlabel metal1 s 0 -48 736 48 8 VGND
port 2 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 3 nsew ground bidirectional
rlabel pwell s 23 21 716 157 6 VNB
port 3 nsew ground bidirectional
rlabel pwell s 532 157 716 203 6 VNB
port 3 nsew ground bidirectional
rlabel nwell s -38 261 774 582 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 496 736 592 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 642 51 719 165 6 X
port 6 nsew signal output
rlabel locali s 663 165 719 299 6 X
port 6 nsew signal output
rlabel locali s 642 299 719 493 6 X
port 6 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 736 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2969424
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2963504
<< end >>
