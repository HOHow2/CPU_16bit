magic
tech sky130A
magscale 1 2
timestamp 1738263620
<< nwell >>
rect -38 261 2246 582
<< pwell >>
rect 1 21 2203 203
rect 30 -17 64 21
<< locali >>
rect 859 323 925 493
rect 1027 323 1093 493
rect 1195 323 1261 493
rect 1363 323 1429 493
rect 1531 323 1597 493
rect 1699 323 1765 493
rect 1867 323 1933 493
rect 2035 323 2101 493
rect 859 289 2191 323
rect 18 215 253 255
rect 2136 181 2191 289
rect 859 147 2191 181
rect 859 52 925 147
rect 859 51 909 52
rect 1027 52 1093 147
rect 1043 51 1077 52
rect 1195 52 1261 147
rect 1211 51 1245 52
rect 1363 52 1429 147
rect 1531 52 1597 147
rect 1699 52 1765 147
rect 1867 52 1933 147
rect 2035 52 2101 147
<< obsli1 >>
rect 0 527 2208 561
rect 19 323 85 493
rect 119 357 153 527
rect 187 323 253 493
rect 287 357 321 527
rect 355 323 421 493
rect 455 367 489 527
rect 523 323 589 493
rect 623 367 657 527
rect 691 323 757 493
rect 791 367 825 527
rect 959 367 993 527
rect 1127 367 1161 527
rect 1295 367 1329 527
rect 1463 367 1497 527
rect 1631 367 1665 527
rect 1799 367 1833 527
rect 1967 367 2001 527
rect 2135 367 2169 527
rect 19 289 321 323
rect 355 289 825 323
rect 287 255 321 289
rect 790 255 825 289
rect 287 215 749 255
rect 790 215 2102 255
rect 287 181 321 215
rect 790 181 825 215
rect 19 147 321 181
rect 355 147 825 181
rect 19 52 85 147
rect 119 17 153 113
rect 187 52 253 147
rect 287 17 321 113
rect 355 52 421 147
rect 455 17 489 113
rect 523 52 589 147
rect 623 17 657 113
rect 691 52 757 147
rect 791 17 825 113
rect 959 17 993 113
rect 1127 17 1161 113
rect 1295 17 1329 113
rect 1463 17 1497 113
rect 1631 17 1665 113
rect 1799 17 1833 113
rect 1967 17 2001 113
rect 2135 17 2169 113
rect 0 -17 2208 17
<< metal1 >>
rect 0 496 2208 592
rect 0 -48 2208 48
<< labels >>
rlabel locali s 18 215 253 255 6 A
port 1 nsew signal input
rlabel metal1 s 0 -48 2208 48 8 VGND
port 2 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 3 nsew ground bidirectional
rlabel pwell s 1 21 2203 203 6 VNB
port 3 nsew ground bidirectional
rlabel nwell s -38 261 2246 582 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 496 2208 592 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 1211 51 1245 52 6 Y
port 6 nsew signal output
rlabel locali s 1043 51 1077 52 6 Y
port 6 nsew signal output
rlabel locali s 859 51 909 52 6 Y
port 6 nsew signal output
rlabel locali s 2035 52 2101 147 6 Y
port 6 nsew signal output
rlabel locali s 1867 52 1933 147 6 Y
port 6 nsew signal output
rlabel locali s 1699 52 1765 147 6 Y
port 6 nsew signal output
rlabel locali s 1531 52 1597 147 6 Y
port 6 nsew signal output
rlabel locali s 1363 52 1429 147 6 Y
port 6 nsew signal output
rlabel locali s 1195 52 1261 147 6 Y
port 6 nsew signal output
rlabel locali s 1027 52 1093 147 6 Y
port 6 nsew signal output
rlabel locali s 859 52 925 147 6 Y
port 6 nsew signal output
rlabel locali s 859 147 2191 181 6 Y
port 6 nsew signal output
rlabel locali s 2136 181 2191 289 6 Y
port 6 nsew signal output
rlabel locali s 859 289 2191 323 6 Y
port 6 nsew signal output
rlabel locali s 2035 323 2101 493 6 Y
port 6 nsew signal output
rlabel locali s 1867 323 1933 493 6 Y
port 6 nsew signal output
rlabel locali s 1699 323 1765 493 6 Y
port 6 nsew signal output
rlabel locali s 1531 323 1597 493 6 Y
port 6 nsew signal output
rlabel locali s 1363 323 1429 493 6 Y
port 6 nsew signal output
rlabel locali s 1195 323 1261 493 6 Y
port 6 nsew signal output
rlabel locali s 1027 323 1093 493 6 Y
port 6 nsew signal output
rlabel locali s 859 323 925 493 6 Y
port 6 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2208 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3280158
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3263332
<< end >>
