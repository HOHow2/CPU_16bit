magic
tech sky130A
magscale 1 2
timestamp 1738263620
<< nwell >>
rect -38 261 1602 582
<< pwell >>
rect 833 157 1563 203
rect 1 21 1563 157
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 351 47 381 131
rect 435 47 465 131
rect 530 47 560 119
rect 628 47 658 119
rect 723 47 753 131
rect 911 47 941 177
rect 1000 47 1030 177
rect 1172 47 1202 177
rect 1360 47 1390 131
rect 1455 47 1485 177
<< scpmoshvt >>
rect 79 363 109 491
rect 163 363 193 491
rect 351 369 381 497
rect 435 369 465 497
rect 531 413 561 497
rect 615 413 645 497
rect 711 413 741 497
rect 908 297 938 497
rect 1000 297 1030 497
rect 1172 297 1202 497
rect 1360 369 1390 497
rect 1455 297 1485 497
<< ndiff >>
rect 27 119 79 131
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 93 163 131
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 119 245 131
rect 193 85 203 119
rect 237 85 245 119
rect 193 47 245 85
rect 299 119 351 131
rect 299 85 307 119
rect 341 85 351 119
rect 299 47 351 85
rect 381 89 435 131
rect 381 55 391 89
rect 425 55 435 89
rect 381 47 435 55
rect 465 119 515 131
rect 673 119 723 131
rect 465 47 530 119
rect 560 107 628 119
rect 560 73 570 107
rect 604 73 628 107
rect 560 47 628 73
rect 658 47 723 119
rect 753 106 805 131
rect 753 72 763 106
rect 797 72 805 106
rect 753 47 805 72
rect 859 129 911 177
rect 859 95 867 129
rect 901 95 911 129
rect 859 47 911 95
rect 941 47 1000 177
rect 1030 89 1172 177
rect 1030 55 1040 89
rect 1074 55 1128 89
rect 1162 55 1172 89
rect 1030 47 1172 55
rect 1202 119 1254 177
rect 1405 131 1455 177
rect 1202 85 1212 119
rect 1246 85 1254 119
rect 1202 47 1254 85
rect 1308 119 1360 131
rect 1308 85 1316 119
rect 1350 85 1360 119
rect 1308 47 1360 85
rect 1390 93 1455 131
rect 1390 59 1411 93
rect 1445 59 1455 93
rect 1390 47 1455 59
rect 1485 103 1537 177
rect 1485 69 1495 103
rect 1529 69 1537 103
rect 1485 47 1537 69
<< pdiff >>
rect 27 477 79 491
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 363 79 375
rect 109 461 163 491
rect 109 427 119 461
rect 153 427 163 461
rect 109 363 163 427
rect 193 477 245 491
rect 193 443 203 477
rect 237 443 245 477
rect 193 409 245 443
rect 193 375 203 409
rect 237 375 245 409
rect 193 363 245 375
rect 299 483 351 497
rect 299 449 307 483
rect 341 449 351 483
rect 299 415 351 449
rect 299 381 307 415
rect 341 381 351 415
rect 299 369 351 381
rect 381 485 435 497
rect 381 451 391 485
rect 425 451 435 485
rect 381 417 435 451
rect 381 383 391 417
rect 425 383 435 417
rect 381 369 435 383
rect 465 413 531 497
rect 561 485 615 497
rect 561 451 571 485
rect 605 451 615 485
rect 561 413 615 451
rect 645 413 711 497
rect 741 477 793 497
rect 741 443 751 477
rect 785 443 793 477
rect 741 413 793 443
rect 856 485 908 497
rect 856 451 864 485
rect 898 451 908 485
rect 465 369 515 413
rect 856 297 908 451
rect 938 471 1000 497
rect 938 437 956 471
rect 990 437 1000 471
rect 938 368 1000 437
rect 938 334 956 368
rect 990 334 1000 368
rect 938 297 1000 334
rect 1030 489 1172 497
rect 1030 455 1040 489
rect 1074 455 1128 489
rect 1162 455 1172 489
rect 1030 421 1172 455
rect 1030 387 1040 421
rect 1074 387 1128 421
rect 1162 387 1172 421
rect 1030 297 1172 387
rect 1202 477 1254 497
rect 1202 443 1212 477
rect 1246 443 1254 477
rect 1202 409 1254 443
rect 1202 375 1212 409
rect 1246 375 1254 409
rect 1202 297 1254 375
rect 1308 450 1360 497
rect 1308 416 1316 450
rect 1350 416 1360 450
rect 1308 369 1360 416
rect 1390 485 1455 497
rect 1390 451 1411 485
rect 1445 451 1455 485
rect 1390 417 1455 451
rect 1390 383 1411 417
rect 1445 383 1455 417
rect 1390 369 1455 383
rect 1405 297 1455 369
rect 1485 477 1537 497
rect 1485 443 1495 477
rect 1529 443 1537 477
rect 1485 409 1537 443
rect 1485 375 1495 409
rect 1529 375 1537 409
rect 1485 297 1537 375
<< ndiffc >>
rect 35 85 69 119
rect 119 59 153 93
rect 203 85 237 119
rect 307 85 341 119
rect 391 55 425 89
rect 570 73 604 107
rect 763 72 797 106
rect 867 95 901 129
rect 1040 55 1074 89
rect 1128 55 1162 89
rect 1212 85 1246 119
rect 1316 85 1350 119
rect 1411 59 1445 93
rect 1495 69 1529 103
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 119 427 153 461
rect 203 443 237 477
rect 203 375 237 409
rect 307 449 341 483
rect 307 381 341 415
rect 391 451 425 485
rect 391 383 425 417
rect 571 451 605 485
rect 751 443 785 477
rect 864 451 898 485
rect 956 437 990 471
rect 956 334 990 368
rect 1040 455 1074 489
rect 1128 455 1162 489
rect 1040 387 1074 421
rect 1128 387 1162 421
rect 1212 443 1246 477
rect 1212 375 1246 409
rect 1316 416 1350 450
rect 1411 451 1445 485
rect 1411 383 1445 417
rect 1495 443 1529 477
rect 1495 375 1529 409
<< poly >>
rect 79 491 109 517
rect 163 491 193 517
rect 351 497 381 523
rect 435 497 465 523
rect 531 497 561 523
rect 615 497 645 523
rect 711 497 741 523
rect 908 497 938 523
rect 1000 497 1030 523
rect 1172 497 1202 523
rect 1360 497 1390 523
rect 1455 497 1485 523
rect 79 348 109 363
rect 45 318 109 348
rect 45 280 75 318
rect 21 264 75 280
rect 163 274 193 363
rect 21 230 31 264
rect 65 230 75 264
rect 21 214 75 230
rect 118 264 193 274
rect 118 230 134 264
rect 168 230 193 264
rect 351 241 381 369
rect 118 220 193 230
rect 45 176 75 214
rect 45 146 109 176
rect 79 131 109 146
rect 163 131 193 220
rect 298 225 381 241
rect 298 191 308 225
rect 342 191 381 225
rect 435 219 465 369
rect 531 337 561 413
rect 615 375 645 413
rect 507 321 561 337
rect 603 365 669 375
rect 603 331 619 365
rect 653 331 669 365
rect 603 321 669 331
rect 711 373 741 413
rect 711 357 812 373
rect 711 323 768 357
rect 802 323 812 357
rect 507 287 517 321
rect 551 287 561 321
rect 711 307 812 323
rect 507 279 561 287
rect 507 271 658 279
rect 531 249 658 271
rect 298 175 381 191
rect 351 131 381 175
rect 424 203 478 219
rect 424 169 434 203
rect 468 169 478 203
rect 424 153 478 169
rect 520 197 586 207
rect 520 163 536 197
rect 570 163 586 197
rect 520 153 586 163
rect 435 131 465 153
rect 530 141 586 153
rect 530 119 560 141
rect 628 119 658 249
rect 723 131 753 307
rect 908 265 938 297
rect 1000 265 1030 297
rect 1172 265 1202 297
rect 1360 265 1390 369
rect 1455 265 1485 297
rect 796 249 941 265
rect 796 215 806 249
rect 840 215 941 249
rect 796 199 941 215
rect 983 249 1037 265
rect 983 215 993 249
rect 1027 215 1037 249
rect 983 199 1037 215
rect 1131 249 1390 265
rect 1131 215 1144 249
rect 1178 215 1390 249
rect 1131 199 1390 215
rect 1435 249 1495 265
rect 1435 215 1445 249
rect 1479 215 1495 249
rect 1435 199 1495 215
rect 911 177 941 199
rect 1000 177 1030 199
rect 1172 177 1202 199
rect 1360 131 1390 199
rect 1455 177 1485 199
rect 79 21 109 47
rect 163 21 193 47
rect 351 21 381 47
rect 435 21 465 47
rect 530 21 560 47
rect 628 21 658 47
rect 723 21 753 47
rect 911 21 941 47
rect 1000 21 1030 47
rect 1172 21 1202 47
rect 1360 21 1390 47
rect 1455 21 1485 47
<< polycont >>
rect 31 230 65 264
rect 134 230 168 264
rect 308 191 342 225
rect 619 331 653 365
rect 768 323 802 357
rect 517 287 551 321
rect 434 169 468 203
rect 536 163 570 197
rect 806 215 840 249
rect 993 215 1027 249
rect 1144 215 1178 249
rect 1445 215 1479 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 17 477 69 493
rect 17 443 35 477
rect 17 409 69 443
rect 103 461 169 527
rect 103 427 119 461
rect 153 427 169 461
rect 203 477 248 493
rect 391 485 454 527
rect 751 485 918 527
rect 1024 489 1178 527
rect 237 443 248 477
rect 17 375 35 409
rect 203 409 248 443
rect 69 375 156 393
rect 17 359 156 375
rect 17 264 65 325
rect 17 230 31 264
rect 17 197 65 230
rect 122 323 156 359
rect 122 280 156 289
rect 237 391 248 409
rect 203 357 214 375
rect 203 337 248 357
rect 291 449 307 483
rect 341 449 357 483
rect 291 415 357 449
rect 291 381 307 415
rect 341 381 357 415
rect 122 264 168 280
rect 122 230 134 264
rect 122 214 168 230
rect 122 161 156 214
rect 17 127 156 161
rect 17 119 69 127
rect 17 85 35 119
rect 203 119 237 337
rect 291 333 357 381
rect 425 451 454 485
rect 549 451 571 485
rect 605 451 717 485
rect 391 417 454 451
rect 654 425 717 451
rect 751 477 864 485
rect 785 451 864 477
rect 898 451 918 485
rect 785 443 918 451
rect 751 427 918 443
rect 956 471 990 487
rect 425 383 454 417
rect 661 415 717 425
rect 679 409 717 415
rect 679 403 721 409
rect 391 367 454 383
rect 585 391 626 399
rect 683 398 721 403
rect 684 395 721 398
rect 686 392 721 395
rect 619 381 626 391
rect 619 365 653 381
rect 291 299 428 333
rect 292 225 358 265
rect 292 191 308 225
rect 342 191 358 225
rect 394 219 428 299
rect 494 323 551 337
rect 528 321 551 323
rect 494 287 517 289
rect 494 271 551 287
rect 585 331 619 357
rect 585 315 653 331
rect 394 203 468 219
rect 585 207 619 315
rect 687 265 721 392
rect 956 373 990 437
rect 1024 455 1040 489
rect 1074 455 1128 489
rect 1162 455 1178 489
rect 1024 421 1178 455
rect 1024 387 1040 421
rect 1074 387 1128 421
rect 1162 387 1178 421
rect 1212 477 1282 493
rect 1246 443 1282 477
rect 1212 409 1282 443
rect 768 368 990 373
rect 768 357 956 368
rect 802 334 956 357
rect 1246 375 1282 409
rect 990 334 1178 353
rect 802 323 1178 334
rect 768 307 1178 323
rect 687 249 840 265
rect 687 233 806 249
rect 394 169 434 203
rect 394 157 468 169
rect 17 69 69 85
rect 103 59 119 93
rect 153 59 169 93
rect 203 69 237 85
rect 307 153 468 157
rect 520 197 619 207
rect 520 163 536 197
rect 570 163 619 197
rect 520 153 619 163
rect 666 215 806 233
rect 666 199 840 215
rect 890 249 1087 265
rect 890 215 993 249
rect 1027 215 1087 249
rect 890 199 1087 215
rect 1131 249 1178 307
rect 1131 215 1144 249
rect 307 123 428 153
rect 307 119 341 123
rect 666 107 700 199
rect 1131 165 1178 215
rect 307 69 341 85
rect 103 17 169 59
rect 375 55 391 89
rect 425 55 441 89
rect 554 73 570 107
rect 604 73 700 107
rect 848 131 1178 165
rect 848 129 908 131
rect 375 17 441 55
rect 747 72 763 106
rect 797 72 814 106
rect 747 17 814 72
rect 848 95 867 129
rect 901 95 908 129
rect 1212 119 1282 375
rect 848 51 908 95
rect 1024 89 1178 97
rect 1024 55 1040 89
rect 1074 55 1128 89
rect 1162 55 1178 89
rect 1024 17 1178 55
rect 1246 85 1282 119
rect 1212 51 1282 85
rect 1316 450 1366 493
rect 1350 416 1366 450
rect 1316 265 1366 416
rect 1402 485 1461 527
rect 1402 451 1411 485
rect 1445 451 1461 485
rect 1402 417 1461 451
rect 1402 383 1411 417
rect 1445 383 1461 417
rect 1402 367 1461 383
rect 1495 477 1547 493
rect 1529 443 1547 477
rect 1495 409 1547 443
rect 1529 375 1547 409
rect 1495 357 1547 375
rect 1316 249 1479 265
rect 1316 215 1445 249
rect 1316 199 1479 215
rect 1316 119 1361 199
rect 1513 119 1547 357
rect 1350 85 1361 119
rect 1495 103 1547 119
rect 1316 51 1361 85
rect 1395 59 1411 93
rect 1445 59 1461 93
rect 1395 17 1461 59
rect 1529 69 1547 103
rect 1495 51 1547 69
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 122 289 156 323
rect 214 375 237 391
rect 237 375 248 391
rect 214 357 248 375
rect 585 357 619 391
rect 494 321 528 323
rect 494 289 517 321
rect 517 289 528 321
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
<< metal1 >>
rect 0 561 1564 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 0 496 1564 527
rect 202 391 260 397
rect 202 357 214 391
rect 248 388 260 391
rect 573 391 631 397
rect 573 388 585 391
rect 248 360 585 388
rect 248 357 260 360
rect 202 351 260 357
rect 573 357 585 360
rect 619 357 631 391
rect 573 351 631 357
rect 110 323 168 329
rect 110 289 122 323
rect 156 320 168 323
rect 482 323 540 329
rect 482 320 494 323
rect 156 292 494 320
rect 156 289 168 292
rect 110 283 168 289
rect 482 289 494 292
rect 528 289 540 323
rect 482 283 540 289
rect 0 17 1564 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
rect 0 -48 1564 -17
<< labels >>
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 GATE
port 2 nsew clock input
flabel locali s 954 221 988 255 0 FreeSans 200 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1500 85 1534 119 0 FreeSans 200 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1046 221 1080 255 0 FreeSans 200 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1220 289 1254 323 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 1220 357 1254 391 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 1220 425 1254 459 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 1220 85 1254 119 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 1500 357 1534 391 0 FreeSans 200 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1220 221 1254 255 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 1500 425 1534 459 0 FreeSans 200 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 310 221 344 255 0 FreeSans 200 0 0 0 D
port 1 nsew signal input
flabel locali s 29 289 63 323 0 FreeSans 200 0 0 0 GATE
port 2 nsew clock input
flabel locali s 1220 153 1254 187 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel nwell s 47 544 47 544 0 FreeSans 200 0 0 0 VPB
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel pwell s 47 0 47 0 0 FreeSans 200 0 0 0 VNB
rlabel comment s 0 0 0 0 4 dlrbp_1
rlabel metal1 s 0 -48 1564 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1564 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1564 544
string GDS_END 2785204
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2771980
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 39.100 0.000 
<< end >>
