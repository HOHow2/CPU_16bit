magic
tech sky130A
magscale 1 2
timestamp 1738263620
<< nwell >>
rect -38 261 2154 582
<< pwell >>
rect 273 157 457 201
rect 1572 181 2041 203
rect 1386 157 2041 181
rect 1 21 2041 157
rect 29 -17 63 21
<< locali >>
rect 18 195 88 325
rect 354 201 436 325
rect 1674 51 1740 493
rect 1973 289 2025 493
rect 1982 165 2025 289
rect 1973 51 2025 165
<< obsli1 >>
rect 0 527 2116 561
rect 35 393 69 493
rect 103 427 169 527
rect 35 359 168 393
rect 122 161 168 359
rect 35 127 168 161
rect 35 69 69 127
rect 103 17 169 93
rect 203 69 248 493
rect 291 427 357 527
rect 391 393 425 493
rect 472 450 638 484
rect 686 451 762 527
rect 286 359 425 393
rect 286 165 320 359
rect 470 315 570 391
rect 286 127 425 165
rect 470 141 514 315
rect 604 281 638 450
rect 798 417 832 475
rect 866 451 932 527
rect 1022 433 1152 483
rect 1186 451 1268 527
rect 1118 417 1152 433
rect 1308 417 1356 475
rect 672 367 942 417
rect 672 315 722 367
rect 824 281 874 313
rect 604 247 874 281
rect 604 239 688 247
rect 550 129 620 203
rect 291 17 357 93
rect 391 61 425 127
rect 654 93 688 239
rect 908 213 942 367
rect 722 147 804 213
rect 862 145 942 213
rect 980 331 1080 393
rect 1118 383 1356 417
rect 1402 389 1468 527
rect 980 179 1014 331
rect 1048 213 1084 295
rect 1118 281 1152 383
rect 1502 353 1536 475
rect 1502 349 1566 353
rect 1186 315 1566 349
rect 1118 247 1494 281
rect 1164 179 1230 203
rect 980 145 1230 179
rect 485 53 688 93
rect 722 17 804 105
rect 862 59 912 145
rect 948 17 1016 109
rect 1264 95 1298 247
rect 1428 235 1494 247
rect 1332 201 1398 213
rect 1332 147 1464 201
rect 1528 136 1566 315
rect 1604 296 1640 527
rect 1128 61 1298 95
rect 1334 17 1466 113
rect 1502 70 1566 136
rect 1604 17 1640 181
rect 1778 265 1844 493
rect 1889 365 1923 527
rect 1778 199 1948 265
rect 1778 51 1844 199
rect 1889 17 1923 117
rect 0 -17 2116 17
<< metal1 >>
rect 0 496 2116 592
rect 753 184 811 193
rect 1397 184 1455 193
rect 753 156 1455 184
rect 753 147 811 156
rect 1397 147 1455 156
rect 0 -48 2116 48
<< obsm1 >>
rect 117 388 175 397
rect 477 388 535 397
rect 1029 388 1087 397
rect 117 360 1087 388
rect 117 351 175 360
rect 477 351 535 360
rect 1029 351 1087 360
rect 1037 252 1095 261
rect 584 224 1095 252
rect 584 193 627 224
rect 1037 215 1095 224
rect 201 184 259 193
rect 569 184 627 193
rect 201 156 627 184
rect 201 147 259 156
rect 569 147 627 156
<< labels >>
rlabel locali s 18 195 88 325 6 CLK
port 1 nsew clock input
rlabel locali s 354 201 436 325 6 D
port 2 nsew signal input
rlabel metal1 s 1397 147 1455 156 6 SET_B
port 3 nsew signal input
rlabel metal1 s 753 147 811 156 6 SET_B
port 3 nsew signal input
rlabel metal1 s 753 156 1455 184 6 SET_B
port 3 nsew signal input
rlabel metal1 s 1397 184 1455 193 6 SET_B
port 3 nsew signal input
rlabel metal1 s 753 184 811 193 6 SET_B
port 3 nsew signal input
rlabel metal1 s 0 -48 2116 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 21 2041 157 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1386 157 2041 181 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1572 181 2041 203 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 273 157 457 201 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 2154 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 2116 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1973 51 2025 165 6 Q
port 8 nsew signal output
rlabel locali s 1982 165 2025 289 6 Q
port 8 nsew signal output
rlabel locali s 1973 289 2025 493 6 Q
port 8 nsew signal output
rlabel locali s 1674 51 1740 493 6 Q_N
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2116 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2571612
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2553846
<< end >>
