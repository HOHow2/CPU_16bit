magic
tech sky130A
magscale 1 2
timestamp 1738263620
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 1 21 624 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 264 47 294 177
rect 348 47 378 177
rect 432 47 462 177
rect 516 47 546 177
<< scpmoshvt >>
rect 91 297 121 497
rect 163 297 193 497
rect 264 297 294 497
rect 348 297 378 497
rect 432 297 462 497
rect 516 297 546 497
<< ndiff >>
rect 27 99 79 177
rect 27 65 35 99
rect 69 65 79 99
rect 27 47 79 65
rect 109 165 163 177
rect 109 131 119 165
rect 153 131 163 165
rect 109 97 163 131
rect 109 63 119 97
rect 153 63 163 97
rect 109 47 163 63
rect 193 132 264 177
rect 193 98 212 132
rect 246 98 264 132
rect 193 47 264 98
rect 294 165 348 177
rect 294 131 304 165
rect 338 131 348 165
rect 294 97 348 131
rect 294 63 304 97
rect 338 63 348 97
rect 294 47 348 63
rect 378 97 432 177
rect 378 63 388 97
rect 422 63 432 97
rect 378 47 432 63
rect 462 165 516 177
rect 462 131 472 165
rect 506 131 516 165
rect 462 97 516 131
rect 462 63 472 97
rect 506 63 516 97
rect 462 47 516 63
rect 546 97 598 177
rect 546 63 556 97
rect 590 63 598 97
rect 546 47 598 63
<< pdiff >>
rect 35 477 91 497
rect 35 443 47 477
rect 81 443 91 477
rect 35 409 91 443
rect 35 375 47 409
rect 81 375 91 409
rect 35 341 91 375
rect 35 307 47 341
rect 81 307 91 341
rect 35 297 91 307
rect 121 297 163 497
rect 193 487 264 497
rect 193 453 212 487
rect 246 453 264 487
rect 193 419 264 453
rect 193 385 212 419
rect 246 385 264 419
rect 193 297 264 385
rect 294 485 348 497
rect 294 451 304 485
rect 338 451 348 485
rect 294 417 348 451
rect 294 383 304 417
rect 338 383 348 417
rect 294 297 348 383
rect 378 485 432 497
rect 378 451 388 485
rect 422 451 432 485
rect 378 297 432 451
rect 462 485 516 497
rect 462 451 472 485
rect 506 451 516 485
rect 462 417 516 451
rect 462 383 472 417
rect 506 383 516 417
rect 462 349 516 383
rect 462 315 472 349
rect 506 315 516 349
rect 462 297 516 315
rect 546 485 602 497
rect 546 451 556 485
rect 590 451 602 485
rect 546 417 602 451
rect 546 383 556 417
rect 590 383 602 417
rect 546 297 602 383
<< ndiffc >>
rect 35 65 69 99
rect 119 131 153 165
rect 119 63 153 97
rect 212 98 246 132
rect 304 131 338 165
rect 304 63 338 97
rect 388 63 422 97
rect 472 131 506 165
rect 472 63 506 97
rect 556 63 590 97
<< pdiffc >>
rect 47 443 81 477
rect 47 375 81 409
rect 47 307 81 341
rect 212 453 246 487
rect 212 385 246 419
rect 304 451 338 485
rect 304 383 338 417
rect 388 451 422 485
rect 472 451 506 485
rect 472 383 506 417
rect 472 315 506 349
rect 556 451 590 485
rect 556 383 590 417
<< poly >>
rect 91 497 121 523
rect 163 497 193 523
rect 264 497 294 523
rect 348 497 378 523
rect 432 497 462 523
rect 516 497 546 523
rect 91 265 121 297
rect 25 249 121 265
rect 25 215 35 249
rect 69 215 121 249
rect 25 199 121 215
rect 163 265 193 297
rect 264 265 294 297
rect 348 265 378 297
rect 432 265 462 297
rect 516 265 546 297
rect 163 249 217 265
rect 163 215 173 249
rect 207 215 217 249
rect 163 199 217 215
rect 264 249 546 265
rect 264 215 298 249
rect 332 215 366 249
rect 400 215 434 249
rect 468 215 546 249
rect 264 199 546 215
rect 79 177 109 199
rect 163 177 193 199
rect 264 177 294 199
rect 348 177 378 199
rect 432 177 462 199
rect 516 177 546 199
rect 79 21 109 47
rect 163 21 193 47
rect 264 21 294 47
rect 348 21 378 47
rect 432 21 462 47
rect 516 21 546 47
<< polycont >>
rect 35 215 69 249
rect 173 215 207 249
rect 298 215 332 249
rect 366 215 400 249
rect 434 215 468 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 31 477 103 493
rect 31 443 47 477
rect 81 443 103 477
rect 31 409 103 443
rect 31 375 47 409
rect 81 375 103 409
rect 31 341 103 375
rect 212 487 246 527
rect 212 419 246 453
rect 212 367 246 385
rect 288 485 354 493
rect 288 451 304 485
rect 338 451 354 485
rect 288 417 354 451
rect 388 485 422 527
rect 388 435 422 451
rect 456 485 522 493
rect 456 451 472 485
rect 506 451 522 485
rect 288 383 304 417
rect 338 401 354 417
rect 456 417 522 451
rect 456 401 472 417
rect 338 383 472 401
rect 506 383 522 417
rect 288 367 522 383
rect 556 485 590 527
rect 556 417 590 451
rect 556 367 590 383
rect 31 307 47 341
rect 81 333 103 341
rect 456 349 522 367
rect 81 307 323 333
rect 31 299 323 307
rect 456 315 472 349
rect 506 333 522 349
rect 506 315 627 333
rect 456 299 627 315
rect 18 249 69 265
rect 18 215 35 249
rect 18 153 69 215
rect 103 165 139 299
rect 173 249 248 265
rect 207 215 248 249
rect 282 249 323 299
rect 282 215 298 249
rect 332 215 366 249
rect 400 215 434 249
rect 468 215 524 249
rect 173 199 248 215
rect 558 181 627 299
rect 288 165 627 181
rect 103 131 119 165
rect 153 131 169 165
rect 21 99 69 119
rect 21 65 35 99
rect 21 17 69 65
rect 103 97 169 131
rect 103 63 119 97
rect 153 63 169 97
rect 103 58 169 63
rect 212 132 246 165
rect 212 17 246 98
rect 288 131 304 165
rect 338 147 472 165
rect 338 131 354 147
rect 288 97 354 131
rect 456 131 472 147
rect 506 147 627 165
rect 506 131 522 147
rect 288 63 304 97
rect 338 63 354 97
rect 288 53 354 63
rect 388 97 422 113
rect 388 17 422 63
rect 456 97 522 131
rect 456 63 472 97
rect 506 63 522 97
rect 456 53 522 63
rect 556 97 590 113
rect 556 17 590 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
flabel locali s 582 289 616 323 0 FreeSans 200 0 0 0 X
port 7 nsew signal output
flabel locali s 214 221 248 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 or2_4
rlabel metal1 s 0 -48 644 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 644 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 644 544
string GDS_END 1003560
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 997858
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 3.220 0.000 
<< end >>
