magic
tech sky130A
magscale 1 2
timestamp 1738263620
<< nwell >>
rect -38 261 1142 582
<< pwell >>
rect 189 157 1085 203
rect 1 21 1085 157
rect 30 -17 64 21
<< locali >>
rect 18 199 66 323
rect 291 333 357 493
rect 459 333 525 493
rect 721 333 787 493
rect 907 333 973 493
rect 291 289 973 333
rect 310 165 357 289
rect 402 215 620 255
rect 672 215 890 255
rect 924 215 1086 255
rect 291 127 357 165
<< obsli1 >>
rect 0 527 1104 561
rect 18 417 69 493
rect 103 451 257 527
rect 18 383 134 417
rect 100 249 134 383
rect 207 289 257 451
rect 391 367 425 527
rect 559 367 687 527
rect 821 367 873 527
rect 1007 299 1086 527
rect 100 215 276 249
rect 100 161 134 215
rect 18 127 134 161
rect 18 51 69 127
rect 207 93 257 181
rect 391 127 609 181
rect 647 143 1068 181
rect 647 127 891 143
rect 391 93 425 127
rect 831 123 891 127
rect 103 17 169 93
rect 207 51 425 93
rect 459 51 797 93
rect 831 51 883 123
rect 933 17 967 109
rect 1001 51 1068 143
rect 0 -17 1104 17
<< metal1 >>
rect 0 496 1104 592
rect 0 -48 1104 48
<< labels >>
rlabel locali s 18 199 66 323 6 A_N
port 1 nsew signal input
rlabel locali s 402 215 620 255 6 B
port 2 nsew signal input
rlabel locali s 672 215 890 255 6 C
port 3 nsew signal input
rlabel locali s 924 215 1086 255 6 D
port 4 nsew signal input
rlabel metal1 s 0 -48 1104 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 21 1085 157 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 189 157 1085 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 1142 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 1104 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 291 127 357 165 6 Y
port 9 nsew signal output
rlabel locali s 310 165 357 289 6 Y
port 9 nsew signal output
rlabel locali s 291 289 973 333 6 Y
port 9 nsew signal output
rlabel locali s 907 333 973 493 6 Y
port 9 nsew signal output
rlabel locali s 721 333 787 493 6 Y
port 9 nsew signal output
rlabel locali s 459 333 525 493 6 Y
port 9 nsew signal output
rlabel locali s 291 333 357 493 6 Y
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1104 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1966168
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1956112
<< end >>
