magic
tech sky130A
magscale 1 2
timestamp 1738263620
<< nwell >>
rect -38 261 1050 582
<< pwell >>
rect 1 21 964 157
rect 29 -17 63 21
<< locali >>
rect 284 347 336 492
rect 456 347 508 492
rect 628 347 680 492
rect 800 347 852 492
rect 284 299 946 347
rect 17 143 80 265
rect 752 181 946 299
rect 284 147 946 181
rect 284 56 336 147
rect 456 56 508 147
rect 628 56 680 147
rect 800 56 852 147
<< obsli1 >>
rect 0 527 1012 561
rect 19 305 78 527
rect 114 265 164 492
rect 198 305 250 527
rect 370 381 422 527
rect 542 381 594 527
rect 714 381 766 527
rect 886 381 945 527
rect 114 215 718 265
rect 29 17 78 109
rect 114 53 164 215
rect 198 17 250 122
rect 370 17 422 113
rect 542 17 594 113
rect 714 17 766 113
rect 886 17 946 113
rect 0 -17 1012 17
<< metal1 >>
rect 0 496 1012 592
rect 0 -48 1012 48
<< labels >>
rlabel locali s 17 143 80 265 6 A
port 1 nsew signal input
rlabel metal1 s 0 -48 1012 48 8 VGND
port 2 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 3 nsew ground bidirectional
rlabel pwell s 1 21 964 157 6 VNB
port 3 nsew ground bidirectional
rlabel nwell s -38 261 1050 582 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 496 1012 592 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 800 56 852 147 6 X
port 6 nsew signal output
rlabel locali s 628 56 680 147 6 X
port 6 nsew signal output
rlabel locali s 456 56 508 147 6 X
port 6 nsew signal output
rlabel locali s 284 56 336 147 6 X
port 6 nsew signal output
rlabel locali s 284 147 946 181 6 X
port 6 nsew signal output
rlabel locali s 752 181 946 299 6 X
port 6 nsew signal output
rlabel locali s 284 299 946 347 6 X
port 6 nsew signal output
rlabel locali s 800 347 852 492 6 X
port 6 nsew signal output
rlabel locali s 628 347 680 492 6 X
port 6 nsew signal output
rlabel locali s 456 347 508 492 6 X
port 6 nsew signal output
rlabel locali s 284 347 336 492 6 X
port 6 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1012 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3293172
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3285430
<< end >>
