magic
tech sky130A
magscale 1 2
timestamp 1738263620
<< nwell >>
rect -38 261 1694 582
<< pwell >>
rect 2 157 272 203
rect 1353 157 1647 203
rect 2 21 1647 157
rect 29 -17 63 21
<< locali >>
rect 120 390 162 493
rect 113 356 162 390
rect 113 317 147 356
rect 17 283 147 317
rect 465 314 683 348
rect 17 181 74 283
rect 17 147 138 181
rect 104 97 138 147
rect 465 255 499 314
rect 425 221 499 255
rect 649 250 683 314
rect 1134 337 1184 391
rect 859 303 1184 337
rect 859 287 931 303
rect 859 250 893 287
rect 1134 271 1184 303
rect 1479 393 1513 493
rect 1479 359 1529 393
rect 649 193 893 250
rect 1495 317 1529 359
rect 1495 283 1639 317
rect 104 63 170 97
rect 1594 181 1639 283
rect 1495 147 1639 181
rect 1495 97 1545 147
rect 1479 51 1545 97
<< obsli1 >>
rect 0 527 1656 561
rect 36 359 70 527
rect 196 455 262 527
rect 380 416 449 493
rect 261 382 449 416
rect 483 421 517 493
rect 551 455 617 527
rect 651 421 698 493
rect 483 387 698 421
rect 739 383 805 527
rect 839 421 873 493
rect 907 455 973 527
rect 1007 421 1041 493
rect 1097 425 1337 493
rect 1378 455 1444 527
rect 839 387 1041 421
rect 1303 421 1337 425
rect 261 333 295 382
rect 188 320 295 333
rect 181 299 295 320
rect 181 286 222 299
rect 329 289 431 338
rect 181 249 215 286
rect 108 215 215 249
rect 36 17 70 113
rect 181 165 215 215
rect 249 255 301 265
rect 249 199 351 255
rect 537 206 615 272
rect 731 287 814 349
rect 1303 387 1436 421
rect 1230 289 1367 347
rect 1402 328 1436 387
rect 1563 359 1597 527
rect 1402 294 1460 328
rect 944 191 1016 255
rect 1050 191 1187 225
rect 1221 199 1392 255
rect 1426 249 1460 294
rect 1426 215 1560 249
rect 385 165 433 187
rect 181 131 433 165
rect 204 17 270 93
rect 307 51 433 131
rect 483 123 685 157
rect 483 51 517 123
rect 551 17 617 89
rect 651 51 685 123
rect 839 123 1041 157
rect 1084 153 1187 191
rect 1426 165 1460 215
rect 739 17 805 98
rect 839 51 873 123
rect 907 17 973 89
rect 1007 51 1041 123
rect 1276 131 1460 165
rect 1108 101 1142 119
rect 1276 101 1310 131
rect 1108 51 1310 101
rect 1356 17 1422 89
rect 1579 17 1613 113
rect 0 -17 1656 17
<< metal1 >>
rect 0 496 1656 592
rect 385 320 443 329
rect 757 320 815 329
rect 1309 320 1367 329
rect 385 292 1367 320
rect 385 283 443 292
rect 757 283 815 292
rect 1309 283 1367 292
rect 293 252 351 261
rect 569 252 627 261
rect 941 252 999 261
rect 1217 252 1275 261
rect 293 224 1275 252
rect 293 215 351 224
rect 569 215 627 224
rect 941 215 999 224
rect 1217 215 1275 224
rect 0 -48 1656 48
<< obsm1 >>
rect 385 184 443 193
rect 1125 184 1183 193
rect 385 156 1183 184
rect 385 147 443 156
rect 1125 147 1183 156
<< labels >>
rlabel metal1 s 1217 215 1275 224 6 A
port 1 nsew signal input
rlabel metal1 s 941 215 999 224 6 A
port 1 nsew signal input
rlabel metal1 s 569 215 627 224 6 A
port 1 nsew signal input
rlabel metal1 s 293 215 351 224 6 A
port 1 nsew signal input
rlabel metal1 s 293 224 1275 252 6 A
port 1 nsew signal input
rlabel metal1 s 1217 252 1275 261 6 A
port 1 nsew signal input
rlabel metal1 s 941 252 999 261 6 A
port 1 nsew signal input
rlabel metal1 s 569 252 627 261 6 A
port 1 nsew signal input
rlabel metal1 s 293 252 351 261 6 A
port 1 nsew signal input
rlabel metal1 s 1309 283 1367 292 6 B
port 2 nsew signal input
rlabel metal1 s 757 283 815 292 6 B
port 2 nsew signal input
rlabel metal1 s 385 283 443 292 6 B
port 2 nsew signal input
rlabel metal1 s 385 292 1367 320 6 B
port 2 nsew signal input
rlabel metal1 s 1309 320 1367 329 6 B
port 2 nsew signal input
rlabel metal1 s 757 320 815 329 6 B
port 2 nsew signal input
rlabel metal1 s 385 320 443 329 6 B
port 2 nsew signal input
rlabel locali s 649 193 893 250 6 CIN
port 3 nsew signal input
rlabel locali s 1134 271 1184 303 6 CIN
port 3 nsew signal input
rlabel locali s 859 250 893 287 6 CIN
port 3 nsew signal input
rlabel locali s 859 287 931 303 6 CIN
port 3 nsew signal input
rlabel locali s 859 303 1184 337 6 CIN
port 3 nsew signal input
rlabel locali s 649 250 683 314 6 CIN
port 3 nsew signal input
rlabel locali s 425 221 499 255 6 CIN
port 3 nsew signal input
rlabel locali s 465 255 499 314 6 CIN
port 3 nsew signal input
rlabel locali s 1134 337 1184 391 6 CIN
port 3 nsew signal input
rlabel locali s 465 314 683 348 6 CIN
port 3 nsew signal input
rlabel metal1 s 0 -48 1656 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 2 21 1647 157 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1353 157 1647 203 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 2 157 272 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 1694 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 1656 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 104 63 170 97 6 COUT
port 8 nsew signal output
rlabel locali s 104 97 138 147 6 COUT
port 8 nsew signal output
rlabel locali s 17 147 138 181 6 COUT
port 8 nsew signal output
rlabel locali s 17 181 74 283 6 COUT
port 8 nsew signal output
rlabel locali s 17 283 147 317 6 COUT
port 8 nsew signal output
rlabel locali s 113 317 147 356 6 COUT
port 8 nsew signal output
rlabel locali s 113 356 162 390 6 COUT
port 8 nsew signal output
rlabel locali s 120 390 162 493 6 COUT
port 8 nsew signal output
rlabel locali s 1479 51 1545 97 6 SUM
port 9 nsew signal output
rlabel locali s 1495 97 1545 147 6 SUM
port 9 nsew signal output
rlabel locali s 1495 147 1639 181 6 SUM
port 9 nsew signal output
rlabel locali s 1594 181 1639 283 6 SUM
port 9 nsew signal output
rlabel locali s 1495 283 1639 317 6 SUM
port 9 nsew signal output
rlabel locali s 1495 317 1529 359 6 SUM
port 9 nsew signal output
rlabel locali s 1479 359 1529 393 6 SUM
port 9 nsew signal output
rlabel locali s 1479 393 1513 493 6 SUM
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1656 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2150438
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2136840
<< end >>
