magic
tech sky130A
magscale 1 2
timestamp 1738263620
<< nwell >>
rect -38 261 1694 582
<< pwell >>
rect 1 21 1655 203
rect 30 -17 64 21
<< locali >>
rect 19 451 757 485
rect 19 97 64 451
rect 1152 285 1570 319
rect 112 221 248 265
rect 112 199 214 221
rect 391 199 710 265
rect 1152 258 1186 285
rect 769 215 1186 258
rect 19 63 757 97
rect 1536 199 1570 285
<< obsli1 >>
rect 0 527 1656 561
rect 795 451 861 527
rect 963 451 1029 527
rect 1131 451 1197 527
rect 1231 417 1265 493
rect 1299 451 1365 527
rect 1399 417 1433 493
rect 1487 451 1553 527
rect 439 383 1433 417
rect 1231 359 1265 383
rect 1399 359 1433 383
rect 1587 359 1639 493
rect 103 315 1116 349
rect 1346 215 1502 249
rect 271 165 340 187
rect 1230 181 1290 187
rect 103 131 340 165
rect 439 131 1097 165
rect 795 17 861 93
rect 895 51 929 131
rect 963 17 1029 93
rect 1063 51 1097 131
rect 1230 143 1433 181
rect 1131 17 1196 118
rect 1230 51 1265 143
rect 1309 17 1359 109
rect 1399 102 1433 143
rect 1468 165 1502 215
rect 1604 165 1639 359
rect 1468 131 1639 165
rect 1487 17 1553 93
rect 1587 51 1639 131
rect 0 -17 1656 17
<< metal1 >>
rect 0 496 1656 592
rect 0 -48 1656 48
<< obsm1 >>
rect 294 184 352 193
rect 1218 184 1276 193
rect 294 156 1276 184
rect 294 147 352 156
rect 1218 147 1276 156
<< labels >>
rlabel locali s 112 199 214 221 6 A0
port 1 nsew signal input
rlabel locali s 112 221 248 265 6 A0
port 1 nsew signal input
rlabel locali s 391 199 710 265 6 A1
port 2 nsew signal input
rlabel locali s 1536 199 1570 285 6 S
port 3 nsew signal input
rlabel locali s 769 215 1186 258 6 S
port 3 nsew signal input
rlabel locali s 1152 258 1186 285 6 S
port 3 nsew signal input
rlabel locali s 1152 285 1570 319 6 S
port 3 nsew signal input
rlabel metal1 s 0 -48 1656 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 21 1655 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 1694 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 1656 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 19 63 757 97 6 Y
port 8 nsew signal output
rlabel locali s 19 97 64 451 6 Y
port 8 nsew signal output
rlabel locali s 19 451 757 485 6 Y
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1656 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1785616
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1773474
<< end >>
