magic
tech sky130A
magscale 1 2
timestamp 1738263620
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 34 21 1195 203
rect 34 17 63 21
rect 29 -17 63 17
<< locali >>
rect 136 333 202 493
rect 304 333 370 493
rect 472 333 538 493
rect 640 333 706 493
rect 808 333 874 493
rect 976 333 1042 493
rect 17 299 1179 333
rect 17 181 102 299
rect 136 215 1054 265
rect 1109 181 1179 299
rect 17 143 1179 181
rect 136 51 202 143
rect 304 51 370 143
rect 472 51 538 143
rect 640 51 706 143
rect 808 51 874 143
rect 976 51 1042 143
<< obsli1 >>
rect 0 527 1196 561
rect 51 367 102 527
rect 236 367 270 527
rect 404 367 438 527
rect 572 367 606 527
rect 740 367 774 527
rect 908 367 942 527
rect 1111 367 1179 527
rect 51 17 102 109
rect 236 17 270 109
rect 404 17 438 109
rect 572 17 606 109
rect 740 17 774 109
rect 908 17 942 109
rect 1111 17 1179 109
rect 0 -17 1196 17
<< metal1 >>
rect 0 496 1196 592
rect 0 -48 1196 48
<< labels >>
rlabel locali s 136 215 1054 265 6 A
port 1 nsew signal input
rlabel metal1 s 0 -48 1196 48 8 VGND
port 2 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 17 8 VNB
port 3 nsew ground bidirectional
rlabel pwell s 34 17 63 21 6 VNB
port 3 nsew ground bidirectional
rlabel pwell s 34 21 1195 203 6 VNB
port 3 nsew ground bidirectional
rlabel nwell s -38 261 1234 582 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 496 1196 592 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 976 51 1042 143 6 Y
port 6 nsew signal output
rlabel locali s 808 51 874 143 6 Y
port 6 nsew signal output
rlabel locali s 640 51 706 143 6 Y
port 6 nsew signal output
rlabel locali s 472 51 538 143 6 Y
port 6 nsew signal output
rlabel locali s 304 51 370 143 6 Y
port 6 nsew signal output
rlabel locali s 136 51 202 143 6 Y
port 6 nsew signal output
rlabel locali s 17 143 1179 181 6 Y
port 6 nsew signal output
rlabel locali s 1109 181 1179 299 6 Y
port 6 nsew signal output
rlabel locali s 17 181 102 299 6 Y
port 6 nsew signal output
rlabel locali s 17 299 1179 333 6 Y
port 6 nsew signal output
rlabel locali s 976 333 1042 493 6 Y
port 6 nsew signal output
rlabel locali s 808 333 874 493 6 Y
port 6 nsew signal output
rlabel locali s 640 333 706 493 6 Y
port 6 nsew signal output
rlabel locali s 472 333 538 493 6 Y
port 6 nsew signal output
rlabel locali s 304 333 370 493 6 Y
port 6 nsew signal output
rlabel locali s 136 333 202 493 6 Y
port 6 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1196 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2250148
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2239840
<< end >>
