magic
tech sky130A
magscale 1 2
timestamp 1738263620
<< nwell >>
rect -38 261 2246 582
<< pwell >>
rect 1175 157 1357 201
rect 1660 157 2196 203
rect 1 145 825 157
rect 1029 145 2196 157
rect 1 21 2196 145
rect 29 -17 63 21
<< locali >>
rect 19 195 89 325
rect 356 157 390 337
rect 492 271 559 337
rect 617 157 651 223
rect 707 207 805 331
rect 356 123 651 157
rect 495 61 530 123
rect 1857 335 1923 479
rect 2027 335 2093 479
rect 1857 301 2191 335
rect 2131 181 2191 301
rect 1857 147 2191 181
rect 1857 61 1923 147
rect 2027 61 2093 147
<< obsli1 >>
rect 0 527 2208 561
rect 36 393 70 493
rect 104 427 170 527
rect 36 359 169 393
rect 123 194 169 359
rect 123 161 162 194
rect 35 127 162 161
rect 204 143 249 493
rect 35 69 69 127
rect 103 17 169 93
rect 203 69 249 143
rect 287 415 342 489
rect 376 449 442 527
rect 539 449 718 483
rect 287 372 650 415
rect 287 89 321 372
rect 424 225 458 372
rect 616 337 650 372
rect 684 399 718 449
rect 752 433 786 527
rect 843 413 890 488
rect 939 438 1153 472
rect 843 399 877 413
rect 684 365 877 399
rect 616 271 655 337
rect 424 191 493 225
rect 843 173 877 365
rect 685 139 877 173
rect 911 207 959 381
rect 997 331 1085 402
rect 1119 315 1153 438
rect 1187 367 1221 527
rect 1255 427 1305 493
rect 1350 433 1527 467
rect 1119 297 1221 315
rect 1061 263 1221 297
rect 911 141 1027 207
rect 287 55 361 89
rect 395 17 461 89
rect 685 89 719 139
rect 843 107 877 139
rect 1061 107 1095 263
rect 1187 249 1221 263
rect 1129 213 1163 219
rect 1255 213 1289 427
rect 1323 249 1361 393
rect 1395 315 1459 381
rect 1129 153 1289 213
rect 1395 207 1433 315
rect 1493 281 1527 433
rect 1563 427 1624 527
rect 1694 381 1751 491
rect 1561 315 1751 381
rect 1785 325 1821 527
rect 1959 369 1993 527
rect 2127 369 2161 527
rect 564 55 719 89
rect 753 17 793 105
rect 843 73 913 107
rect 947 73 1095 107
rect 1145 17 1219 117
rect 1255 107 1289 153
rect 1323 141 1433 207
rect 1467 265 1527 281
rect 1714 265 1751 315
rect 1467 199 1680 265
rect 1714 215 2097 265
rect 1467 107 1501 199
rect 1714 165 1750 215
rect 1255 73 1347 107
rect 1393 73 1501 107
rect 1550 17 1624 123
rect 1678 60 1750 165
rect 1785 17 1819 139
rect 1959 17 1993 113
rect 2127 17 2161 113
rect 0 -17 2208 17
<< metal1 >>
rect 0 496 2208 592
rect 0 -48 2208 48
<< obsm1 >>
rect 111 388 169 397
rect 1031 388 1089 397
rect 1313 388 1371 397
rect 111 360 1371 388
rect 111 351 169 360
rect 1031 351 1089 360
rect 1313 351 1371 360
rect 199 184 257 193
rect 939 184 997 193
rect 1313 184 1371 193
rect 199 156 1371 184
rect 199 147 257 156
rect 939 147 997 156
rect 1313 147 1371 156
<< labels >>
rlabel locali s 19 195 89 325 6 CLK
port 1 nsew clock input
rlabel locali s 492 271 559 337 6 D
port 2 nsew signal input
rlabel locali s 707 207 805 331 6 SCD
port 3 nsew signal input
rlabel locali s 495 61 530 123 6 SCE
port 4 nsew signal input
rlabel locali s 356 123 651 157 6 SCE
port 4 nsew signal input
rlabel locali s 617 157 651 223 6 SCE
port 4 nsew signal input
rlabel locali s 356 157 390 337 6 SCE
port 4 nsew signal input
rlabel metal1 s 0 -48 2208 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 21 2196 145 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1029 145 2196 157 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 145 825 157 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1660 157 2196 203 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1175 157 1357 201 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 2246 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 2208 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 2027 61 2093 147 6 Q
port 9 nsew signal output
rlabel locali s 1857 61 1923 147 6 Q
port 9 nsew signal output
rlabel locali s 1857 147 2191 181 6 Q
port 9 nsew signal output
rlabel locali s 2131 181 2191 301 6 Q
port 9 nsew signal output
rlabel locali s 1857 301 2191 335 6 Q
port 9 nsew signal output
rlabel locali s 2027 335 2093 479 6 Q
port 9 nsew signal output
rlabel locali s 1857 335 1923 479 6 Q
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2208 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 408676
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 392218
<< end >>
