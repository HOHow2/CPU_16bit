magic
tech sky130A
magscale 1 2
timestamp 1738263620
<< nwell >>
rect -38 261 1694 582
<< pwell >>
rect 834 157 1655 203
rect 1 21 1655 157
rect 30 -17 64 21
<< locali >>
rect 17 197 66 325
rect 292 191 358 265
rect 1136 332 1186 493
rect 1136 299 1213 332
rect 1158 265 1213 299
rect 1503 321 1553 493
rect 1519 265 1553 321
rect 880 199 1030 265
rect 1158 177 1272 265
rect 1519 211 1639 265
rect 1158 167 1230 177
rect 1136 133 1230 167
rect 1136 66 1170 133
rect 1519 165 1553 211
rect 1503 51 1553 165
<< obsli1 >>
rect 0 527 1656 561
rect 17 393 69 493
rect 103 427 169 527
rect 17 359 156 393
rect 122 280 156 359
rect 203 337 248 493
rect 122 214 168 280
rect 122 161 156 214
rect 17 127 156 161
rect 17 69 69 127
rect 103 17 169 93
rect 203 69 237 337
rect 291 333 357 483
rect 391 367 454 527
rect 549 451 717 485
rect 654 425 717 451
rect 751 427 920 527
rect 661 415 717 425
rect 679 409 717 415
rect 679 403 721 409
rect 585 381 625 399
rect 683 398 721 403
rect 684 395 721 398
rect 686 392 721 395
rect 291 299 428 333
rect 394 219 428 299
rect 494 271 551 337
rect 585 315 653 381
rect 394 157 468 219
rect 585 207 619 315
rect 687 265 721 392
rect 954 373 988 487
rect 1022 375 1098 527
rect 768 341 988 373
rect 768 307 1102 341
rect 1064 265 1102 307
rect 1220 366 1272 527
rect 1307 265 1374 493
rect 1409 367 1468 527
rect 1587 299 1639 527
rect 687 233 840 265
rect 307 153 468 157
rect 307 123 428 153
rect 543 141 619 207
rect 666 199 840 233
rect 1064 199 1124 265
rect 307 69 341 123
rect 666 107 700 199
rect 1064 165 1102 199
rect 1307 199 1485 265
rect 375 17 441 89
rect 554 73 700 107
rect 854 131 1102 165
rect 748 17 814 106
rect 854 83 914 131
rect 1022 17 1098 97
rect 1204 17 1272 93
rect 1307 51 1373 199
rect 1407 17 1468 109
rect 1587 17 1639 177
rect 0 -17 1656 17
<< metal1 >>
rect 0 496 1656 592
rect 0 -48 1656 48
<< obsm1 >>
rect 202 388 260 397
rect 574 388 632 397
rect 202 360 632 388
rect 202 351 260 360
rect 574 351 632 360
rect 110 320 168 329
rect 482 320 540 329
rect 110 292 540 320
rect 110 283 168 292
rect 482 283 540 292
<< labels >>
rlabel locali s 292 191 358 265 6 D
port 1 nsew signal input
rlabel locali s 17 197 66 325 6 GATE
port 2 nsew clock input
rlabel locali s 880 199 1030 265 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 0 -48 1656 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 21 1655 157 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 834 157 1655 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 1694 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 1656 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1136 66 1170 133 6 Q
port 8 nsew signal output
rlabel locali s 1136 133 1230 167 6 Q
port 8 nsew signal output
rlabel locali s 1158 167 1230 177 6 Q
port 8 nsew signal output
rlabel locali s 1158 177 1272 265 6 Q
port 8 nsew signal output
rlabel locali s 1158 265 1213 299 6 Q
port 8 nsew signal output
rlabel locali s 1136 299 1213 332 6 Q
port 8 nsew signal output
rlabel locali s 1136 332 1186 493 6 Q
port 8 nsew signal output
rlabel locali s 1503 51 1553 165 6 Q_N
port 9 nsew signal output
rlabel locali s 1519 165 1553 211 6 Q_N
port 9 nsew signal output
rlabel locali s 1519 211 1639 265 6 Q_N
port 9 nsew signal output
rlabel locali s 1519 265 1553 321 6 Q_N
port 9 nsew signal output
rlabel locali s 1503 321 1553 493 6 Q_N
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1656 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2800102
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2785260
<< end >>
