magic
tech sky130A
magscale 1 2
timestamp 1738263620
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 1 67 735 203
rect 29 21 735 67
rect 29 -17 63 21
<< locali >>
rect 119 265 155 339
rect 85 199 155 265
rect 189 299 270 339
rect 189 119 223 299
rect 489 215 586 257
rect 620 215 719 325
rect 189 51 248 119
<< obsli1 >>
rect 0 527 736 561
rect 104 441 182 527
rect 283 441 446 527
rect 480 407 545 493
rect 17 373 387 407
rect 17 299 79 373
rect 17 165 51 299
rect 17 86 69 165
rect 119 17 155 165
rect 257 212 291 265
rect 257 178 319 212
rect 353 199 387 373
rect 421 291 545 407
rect 640 375 706 527
rect 285 165 319 178
rect 421 165 455 291
rect 285 131 455 165
rect 282 17 354 97
rect 388 51 455 131
rect 489 147 718 181
rect 489 73 549 147
rect 583 17 617 111
rect 651 54 718 147
rect 0 -17 736 17
<< metal1 >>
rect 0 496 736 592
rect 0 -48 736 48
<< labels >>
rlabel locali s 620 215 719 325 6 A1
port 1 nsew signal input
rlabel locali s 489 215 586 257 6 A2
port 2 nsew signal input
rlabel locali s 85 199 155 265 6 B1_N
port 3 nsew signal input
rlabel locali s 119 265 155 339 6 B1_N
port 3 nsew signal input
rlabel metal1 s 0 -48 736 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 29 21 735 67 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 67 735 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 774 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 736 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 189 51 248 119 6 X
port 8 nsew signal output
rlabel locali s 189 119 223 299 6 X
port 8 nsew signal output
rlabel locali s 189 299 270 339 6 X
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 736 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1338728
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1332440
<< end >>
