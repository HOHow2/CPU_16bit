magic
tech sky130A
magscale 1 2
timestamp 1738263620
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 1 21 919 203
rect 30 -17 64 21
<< locali >>
rect 751 323 817 423
rect 29 199 164 323
rect 210 199 351 323
rect 391 199 533 323
rect 651 289 817 323
rect 581 199 615 265
rect 651 165 714 289
rect 853 255 898 325
rect 764 215 898 255
rect 459 131 901 165
rect 651 51 685 131
rect 835 59 901 131
<< obsli1 >>
rect 0 527 920 561
rect 35 391 69 493
rect 103 425 169 527
rect 203 391 237 493
rect 271 425 337 527
rect 371 391 405 493
rect 462 425 596 527
rect 667 459 885 493
rect 667 391 701 459
rect 35 357 701 391
rect 851 359 885 459
rect 19 131 421 165
rect 103 17 169 93
rect 271 59 615 93
rect 735 17 801 93
rect 0 -17 920 17
<< metal1 >>
rect 0 496 920 592
rect 0 -48 920 48
<< labels >>
rlabel locali s 581 199 615 265 6 A1
port 1 nsew signal input
rlabel locali s 391 199 533 323 6 A1
port 1 nsew signal input
rlabel locali s 210 199 351 323 6 A2
port 2 nsew signal input
rlabel locali s 29 199 164 323 6 A3
port 3 nsew signal input
rlabel locali s 764 215 898 255 6 B1
port 4 nsew signal input
rlabel locali s 853 255 898 325 6 B1
port 4 nsew signal input
rlabel metal1 s 0 -48 920 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 21 919 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 958 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 920 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 835 59 901 131 6 Y
port 9 nsew signal output
rlabel locali s 651 51 685 131 6 Y
port 9 nsew signal output
rlabel locali s 459 131 901 165 6 Y
port 9 nsew signal output
rlabel locali s 651 165 714 289 6 Y
port 9 nsew signal output
rlabel locali s 651 289 817 323 6 Y
port 9 nsew signal output
rlabel locali s 751 323 817 423 6 Y
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 920 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3503672
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3494670
<< end >>
