magic
tech sky130A
magscale 1 2
timestamp 1738263620
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 1 157 187 203
rect 735 157 919 203
rect 1 21 919 157
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 267 47 297 131
rect 351 47 381 131
rect 435 47 465 131
rect 644 47 674 131
rect 716 47 746 131
rect 811 47 841 177
<< scpmoshvt >>
rect 79 297 109 497
rect 262 413 292 497
rect 346 413 376 497
rect 456 413 486 497
rect 628 413 658 497
rect 716 413 746 497
rect 811 297 841 497
<< ndiff >>
rect 27 165 79 177
rect 27 131 35 165
rect 69 131 79 165
rect 27 97 79 131
rect 27 63 35 97
rect 69 63 79 97
rect 27 47 79 63
rect 109 161 161 177
rect 109 127 119 161
rect 153 127 161 161
rect 761 131 811 177
rect 109 93 161 127
rect 109 59 119 93
rect 153 59 161 93
rect 109 47 161 59
rect 215 119 267 131
rect 215 85 223 119
rect 257 85 267 119
rect 215 47 267 85
rect 297 119 351 131
rect 297 85 307 119
rect 341 85 351 119
rect 297 47 351 85
rect 381 93 435 131
rect 381 59 391 93
rect 425 59 435 93
rect 381 47 435 59
rect 465 119 517 131
rect 465 85 475 119
rect 509 85 517 119
rect 465 47 517 85
rect 592 119 644 131
rect 592 85 600 119
rect 634 85 644 119
rect 592 47 644 85
rect 674 47 716 131
rect 746 93 811 131
rect 746 59 767 93
rect 801 59 811 93
rect 746 47 811 59
rect 841 165 893 177
rect 841 131 851 165
rect 885 131 893 165
rect 841 97 893 131
rect 841 63 851 97
rect 885 63 893 97
rect 841 47 893 63
<< pdiff >>
rect 27 483 79 497
rect 27 449 35 483
rect 69 449 79 483
rect 27 415 79 449
rect 27 381 35 415
rect 69 381 79 415
rect 27 347 79 381
rect 27 313 35 347
rect 69 313 79 347
rect 27 297 79 313
rect 109 489 262 497
rect 109 455 119 489
rect 153 455 202 489
rect 236 455 262 489
rect 109 421 262 455
rect 109 387 119 421
rect 153 413 262 421
rect 292 455 346 497
rect 292 421 302 455
rect 336 421 346 455
rect 292 413 346 421
rect 376 413 456 497
rect 486 489 628 497
rect 486 455 506 489
rect 540 455 574 489
rect 608 455 628 489
rect 486 413 628 455
rect 658 455 716 497
rect 658 421 670 455
rect 704 421 716 455
rect 658 413 716 421
rect 746 475 811 497
rect 746 441 767 475
rect 801 441 811 475
rect 746 413 811 441
rect 153 387 161 413
rect 109 353 161 387
rect 109 319 119 353
rect 153 319 161 353
rect 109 297 161 319
rect 761 297 811 413
rect 841 483 893 497
rect 841 449 851 483
rect 885 449 893 483
rect 841 415 893 449
rect 841 381 851 415
rect 885 381 893 415
rect 841 347 893 381
rect 841 313 851 347
rect 885 313 893 347
rect 841 297 893 313
<< ndiffc >>
rect 35 131 69 165
rect 35 63 69 97
rect 119 127 153 161
rect 119 59 153 93
rect 223 85 257 119
rect 307 85 341 119
rect 391 59 425 93
rect 475 85 509 119
rect 600 85 634 119
rect 767 59 801 93
rect 851 131 885 165
rect 851 63 885 97
<< pdiffc >>
rect 35 449 69 483
rect 35 381 69 415
rect 35 313 69 347
rect 119 455 153 489
rect 202 455 236 489
rect 119 387 153 421
rect 302 421 336 455
rect 506 455 540 489
rect 574 455 608 489
rect 670 421 704 455
rect 767 441 801 475
rect 119 319 153 353
rect 851 449 885 483
rect 851 381 885 415
rect 851 313 885 347
<< poly >>
rect 79 497 109 523
rect 262 497 292 523
rect 346 497 376 523
rect 456 497 486 523
rect 628 497 658 523
rect 716 497 746 523
rect 811 497 841 523
rect 79 265 109 297
rect 262 265 292 413
rect 346 365 376 413
rect 346 349 414 365
rect 346 315 370 349
rect 404 315 414 349
rect 346 299 414 315
rect 456 313 486 413
rect 628 385 658 413
rect 597 381 658 385
rect 573 365 658 381
rect 573 331 583 365
rect 617 355 658 365
rect 617 331 627 355
rect 573 315 627 331
rect 79 249 158 265
rect 79 215 114 249
rect 148 215 158 249
rect 79 199 158 215
rect 250 249 304 265
rect 250 215 260 249
rect 294 215 304 249
rect 250 199 304 215
rect 79 177 109 199
rect 267 131 297 199
rect 351 131 381 299
rect 456 297 527 313
rect 456 263 483 297
rect 517 263 527 297
rect 456 257 527 263
rect 434 247 527 257
rect 434 227 486 247
rect 435 131 465 227
rect 597 177 627 315
rect 716 297 746 413
rect 669 281 746 297
rect 669 247 679 281
rect 713 247 746 281
rect 811 265 841 297
rect 669 231 746 247
rect 597 147 674 177
rect 644 131 674 147
rect 716 131 746 231
rect 788 249 842 265
rect 788 215 798 249
rect 832 215 842 249
rect 788 199 842 215
rect 811 177 841 199
rect 79 21 109 47
rect 267 21 297 47
rect 351 21 381 47
rect 435 21 465 47
rect 644 21 674 47
rect 716 21 746 47
rect 811 21 841 47
<< polycont >>
rect 370 315 404 349
rect 583 331 617 365
rect 114 215 148 249
rect 260 215 294 249
rect 483 263 517 297
rect 679 247 713 281
rect 798 215 832 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 119 489 252 527
rect 18 449 35 483
rect 69 449 85 483
rect 18 415 85 449
rect 18 381 35 415
rect 69 381 85 415
rect 18 347 85 381
rect 18 313 35 347
rect 69 313 85 347
rect 153 455 202 489
rect 236 455 252 489
rect 490 489 624 527
rect 302 455 336 471
rect 119 421 158 455
rect 153 387 158 421
rect 119 353 158 387
rect 153 319 158 353
rect 18 165 64 313
rect 119 303 158 319
rect 192 387 336 421
rect 192 249 226 387
rect 370 365 431 475
rect 490 455 506 489
rect 540 455 574 489
rect 608 455 624 489
rect 751 475 801 527
rect 670 455 704 471
rect 751 441 767 475
rect 751 425 801 441
rect 835 449 851 483
rect 885 449 903 483
rect 670 391 704 421
rect 835 415 903 449
rect 370 349 583 365
rect 404 331 583 349
rect 617 331 633 365
rect 670 357 801 391
rect 404 315 431 331
rect 370 269 431 315
rect 672 297 717 323
rect 98 215 114 249
rect 148 215 226 249
rect 18 131 35 165
rect 69 131 85 165
rect 18 97 85 131
rect 18 63 35 97
rect 69 63 85 97
rect 119 161 158 177
rect 153 127 158 161
rect 119 93 158 127
rect 153 59 158 93
rect 192 135 226 215
rect 260 249 294 265
rect 467 263 483 297
rect 517 281 717 297
rect 517 263 679 281
rect 672 247 679 263
rect 713 247 717 281
rect 294 215 634 229
rect 260 195 634 215
rect 672 211 717 247
rect 767 265 801 357
rect 835 381 851 415
rect 885 381 903 415
rect 835 347 903 381
rect 835 313 851 347
rect 885 313 903 347
rect 767 249 832 265
rect 767 215 798 249
rect 600 177 634 195
rect 767 199 832 215
rect 767 177 801 199
rect 192 119 257 135
rect 192 85 223 119
rect 192 69 257 85
rect 307 127 509 161
rect 307 119 341 127
rect 475 119 509 127
rect 307 69 341 85
rect 119 17 158 59
rect 375 59 391 93
rect 425 59 441 93
rect 475 69 509 85
rect 600 143 801 177
rect 866 165 903 313
rect 600 119 634 143
rect 835 131 851 165
rect 885 131 903 165
rect 600 69 634 85
rect 751 93 801 109
rect 375 17 441 59
rect 751 59 767 93
rect 835 97 903 131
rect 835 63 851 97
rect 885 63 903 97
rect 751 17 801 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel locali s 397 425 431 459 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 672 221 706 255 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 856 357 890 391 0 FreeSans 340 0 0 0 COUT
port 7 nsew signal output
flabel locali s 856 85 890 119 0 FreeSans 340 0 0 0 COUT
port 7 nsew signal output
flabel locali s 30 85 64 119 0 FreeSans 340 0 0 0 SUM
port 8 nsew signal output
flabel locali s 30 153 64 187 0 FreeSans 340 0 0 0 SUM
port 8 nsew signal output
flabel locali s 30 221 64 255 0 FreeSans 340 0 0 0 SUM
port 8 nsew signal output
flabel locali s 30 289 64 323 0 FreeSans 340 0 0 0 SUM
port 8 nsew signal output
flabel locali s 30 357 64 391 0 FreeSans 340 0 0 0 SUM
port 8 nsew signal output
flabel locali s 30 425 64 459 0 FreeSans 340 0 0 0 SUM
port 8 nsew signal output
flabel locali s 856 425 890 459 0 FreeSans 340 0 0 0 COUT
port 7 nsew signal output
flabel locali s 672 289 706 323 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 397 357 431 391 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 397 289 431 323 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
rlabel comment s 0 0 0 0 4 ha_1
rlabel metal1 s 0 -48 920 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 920 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 920 544
string GDS_END 2304928
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2296048
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 12.300 1.725 12.300 3.600 8.100 3.600 8.100 1.725 
<< end >>
