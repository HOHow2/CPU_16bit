magic
tech sky130A
magscale 1 2
timestamp 1738263620
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 3 157 272 203
rect 3 21 808 157
rect 25 -17 59 21
<< locali >>
rect 105 305 156 493
rect 105 162 139 305
rect 269 199 335 323
rect 369 199 427 275
rect 105 51 156 162
rect 610 271 706 331
rect 654 153 706 271
rect 746 153 798 331
<< obsli1 >>
rect 0 527 828 561
rect 37 289 71 527
rect 190 447 256 527
rect 500 474 534 493
rect 308 440 534 474
rect 575 451 641 485
rect 308 395 342 440
rect 190 361 342 395
rect 488 413 534 440
rect 37 17 71 186
rect 190 265 224 361
rect 395 343 429 381
rect 488 379 570 413
rect 173 199 224 265
rect 395 309 502 343
rect 468 165 502 309
rect 323 131 502 165
rect 536 174 570 379
rect 607 401 641 451
rect 675 435 725 527
rect 759 401 793 493
rect 607 367 793 401
rect 536 140 606 174
rect 190 17 276 106
rect 323 51 357 131
rect 391 17 538 97
rect 572 51 606 140
rect 721 17 801 119
rect 0 -17 828 17
<< metal1 >>
rect 0 496 828 592
rect 0 -48 828 48
<< labels >>
rlabel locali s 269 199 335 323 6 A1_N
port 1 nsew signal input
rlabel locali s 369 199 427 275 6 A2_N
port 2 nsew signal input
rlabel locali s 746 153 798 331 6 B1
port 3 nsew signal input
rlabel locali s 654 153 706 271 6 B2
port 4 nsew signal input
rlabel locali s 610 271 706 331 6 B2
port 4 nsew signal input
rlabel metal1 s 0 -48 828 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 25 -17 59 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 3 21 808 157 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 3 157 272 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 866 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 828 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 105 51 156 162 6 X
port 9 nsew signal output
rlabel locali s 105 162 139 305 6 X
port 9 nsew signal output
rlabel locali s 105 305 156 493 6 X
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 828 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3986106
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3978378
<< end >>
