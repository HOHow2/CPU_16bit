magic
tech sky130A
magscale 1 2
timestamp 1738263620
<< nwell >>
rect -38 261 590 582
<< pwell >>
rect 1 21 551 203
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 177
rect 267 47 297 177
rect 359 47 389 177
rect 443 47 473 177
<< scpmoshvt >>
rect 83 297 113 497
rect 244 297 274 497
rect 352 297 382 497
rect 443 297 473 497
<< ndiff >>
rect 27 164 79 177
rect 27 130 35 164
rect 69 130 79 164
rect 27 96 79 130
rect 27 62 35 96
rect 69 62 79 96
rect 27 47 79 62
rect 109 93 161 177
rect 109 59 119 93
rect 153 59 161 93
rect 109 47 161 59
rect 215 165 267 177
rect 215 131 223 165
rect 257 131 267 165
rect 215 97 267 131
rect 215 63 223 97
rect 257 63 267 97
rect 215 47 267 63
rect 297 161 359 177
rect 297 127 315 161
rect 349 127 359 161
rect 297 47 359 127
rect 389 93 443 177
rect 389 59 399 93
rect 433 59 443 93
rect 389 47 443 59
rect 473 165 525 177
rect 473 131 483 165
rect 517 131 525 165
rect 473 97 525 131
rect 473 63 483 97
rect 517 63 525 97
rect 473 47 525 63
<< pdiff >>
rect 27 477 83 497
rect 27 443 39 477
rect 73 443 83 477
rect 27 409 83 443
rect 27 375 39 409
rect 73 375 83 409
rect 27 341 83 375
rect 27 307 39 341
rect 73 307 83 341
rect 27 297 83 307
rect 113 485 244 497
rect 113 451 125 485
rect 159 451 199 485
rect 233 451 244 485
rect 113 417 244 451
rect 113 383 125 417
rect 159 383 199 417
rect 233 383 244 417
rect 113 297 244 383
rect 274 485 352 497
rect 274 451 299 485
rect 333 451 352 485
rect 274 417 352 451
rect 274 383 299 417
rect 333 383 352 417
rect 274 349 352 383
rect 274 315 299 349
rect 333 315 352 349
rect 274 297 352 315
rect 382 297 443 497
rect 473 485 525 497
rect 473 451 483 485
rect 517 451 525 485
rect 473 417 525 451
rect 473 383 483 417
rect 517 383 525 417
rect 473 297 525 383
<< ndiffc >>
rect 35 130 69 164
rect 35 62 69 96
rect 119 59 153 93
rect 223 131 257 165
rect 223 63 257 97
rect 315 127 349 161
rect 399 59 433 93
rect 483 131 517 165
rect 483 63 517 97
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 39 307 73 341
rect 125 451 159 485
rect 199 451 233 485
rect 125 383 159 417
rect 199 383 233 417
rect 299 451 333 485
rect 299 383 333 417
rect 299 315 333 349
rect 483 451 517 485
rect 483 383 517 417
<< poly >>
rect 83 497 113 523
rect 244 497 274 523
rect 352 497 382 523
rect 443 497 473 523
rect 83 265 113 297
rect 244 265 274 297
rect 352 265 382 297
rect 443 269 473 297
rect 79 249 163 265
rect 79 215 119 249
rect 153 215 163 249
rect 79 199 163 215
rect 244 249 301 265
rect 244 215 257 249
rect 291 215 301 249
rect 244 199 301 215
rect 347 249 401 265
rect 347 215 357 249
rect 391 215 401 249
rect 347 199 401 215
rect 443 249 529 269
rect 443 215 485 249
rect 519 215 529 249
rect 443 199 529 215
rect 79 177 109 199
rect 267 177 297 199
rect 359 177 389 199
rect 443 177 473 199
rect 79 21 109 47
rect 267 21 297 47
rect 359 21 389 47
rect 443 21 473 47
<< polycont >>
rect 119 215 153 249
rect 257 215 291 249
rect 357 215 391 249
rect 485 215 519 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 17 477 73 493
rect 17 443 39 477
rect 17 409 73 443
rect 17 375 39 409
rect 17 341 73 375
rect 107 485 249 527
rect 107 451 125 485
rect 159 451 199 485
rect 233 451 249 485
rect 107 417 249 451
rect 107 383 125 417
rect 159 383 199 417
rect 233 383 249 417
rect 107 372 249 383
rect 283 485 349 493
rect 283 451 299 485
rect 333 451 349 485
rect 467 485 533 527
rect 283 417 349 451
rect 283 383 299 417
rect 333 383 349 417
rect 17 307 39 341
rect 283 349 349 383
rect 283 338 299 349
rect 17 206 73 307
rect 119 315 299 338
rect 333 315 349 349
rect 119 295 349 315
rect 119 249 176 295
rect 153 215 176 249
rect 213 249 307 261
rect 388 255 431 478
rect 467 451 483 485
rect 517 451 533 485
rect 467 417 533 451
rect 467 383 483 417
rect 517 383 533 417
rect 489 255 535 323
rect 213 215 257 249
rect 291 215 307 249
rect 341 249 431 255
rect 341 215 357 249
rect 391 219 431 249
rect 469 249 535 255
rect 391 215 407 219
rect 469 215 485 249
rect 519 215 535 249
rect 17 164 85 206
rect 17 130 35 164
rect 69 130 85 164
rect 119 181 176 215
rect 119 165 261 181
rect 119 143 223 165
rect 17 96 85 130
rect 201 131 223 143
rect 257 131 261 165
rect 201 115 261 131
rect 299 165 535 181
rect 299 161 483 165
rect 299 127 315 161
rect 349 143 483 161
rect 349 127 365 143
rect 467 131 483 143
rect 517 131 535 165
rect 201 113 264 115
rect 201 111 266 113
rect 201 110 268 111
rect 17 62 35 96
rect 69 62 85 96
rect 17 51 85 62
rect 119 93 153 109
rect 119 17 153 59
rect 201 108 269 110
rect 201 107 270 108
rect 201 105 271 107
rect 201 104 272 105
rect 201 97 273 104
rect 201 63 223 97
rect 257 63 273 97
rect 201 51 273 63
rect 399 93 433 109
rect 399 17 433 59
rect 467 97 535 131
rect 467 63 483 97
rect 517 63 535 97
rect 467 51 535 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
<< metal1 >>
rect 0 561 552 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 0 496 552 527
rect 0 17 552 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
rect 0 -48 552 -17
<< labels >>
flabel locali s 29 357 63 391 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 489 289 523 323 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 213 221 247 255 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 397 221 431 255 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 o21a_1
rlabel metal1 s 0 -48 552 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 552 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 552 544
string GDS_END 1296620
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1291048
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 2.760 0.000 
<< end >>
