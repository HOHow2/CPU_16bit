* NGSPICE file created from sky130_ef_sc_hd__fill_2.ext - technology: sky130A

.subckt sky130_ef_sc_hd__fill_2 VNB VPB VGND VPWR
.ends

