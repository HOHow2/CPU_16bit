magic
tech sky130A
magscale 1 2
timestamp 1738263620
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 6 21 1152 203
rect 29 -17 63 21
<< scnmos >>
rect 85 47 115 177
rect 171 47 201 177
rect 257 47 287 177
rect 343 47 373 177
rect 429 47 459 177
rect 515 47 545 177
rect 601 47 631 177
rect 695 47 725 177
rect 781 47 811 177
rect 867 47 897 177
rect 953 47 983 177
rect 1039 47 1069 177
<< scpmoshvt >>
rect 85 297 115 497
rect 171 297 201 497
rect 257 297 287 497
rect 343 297 373 497
rect 429 297 459 497
rect 515 297 545 497
rect 601 297 631 497
rect 687 297 717 497
rect 781 297 811 497
rect 867 297 897 497
rect 953 297 983 497
rect 1039 297 1069 497
<< ndiff >>
rect 32 157 85 177
rect 32 123 40 157
rect 74 123 85 157
rect 32 47 85 123
rect 115 89 171 177
rect 115 55 126 89
rect 160 55 171 89
rect 115 47 171 55
rect 201 157 257 177
rect 201 123 212 157
rect 246 123 257 157
rect 201 47 257 123
rect 287 89 343 177
rect 287 55 298 89
rect 332 55 343 89
rect 287 47 343 55
rect 373 157 429 177
rect 373 123 384 157
rect 418 123 429 157
rect 373 47 429 123
rect 459 89 515 177
rect 459 55 470 89
rect 504 55 515 89
rect 459 47 515 55
rect 545 157 601 177
rect 545 123 556 157
rect 590 123 601 157
rect 545 47 601 123
rect 631 89 695 177
rect 631 55 642 89
rect 676 55 695 89
rect 631 47 695 55
rect 725 125 781 177
rect 725 91 736 125
rect 770 91 781 125
rect 725 47 781 91
rect 811 157 867 177
rect 811 123 822 157
rect 856 123 867 157
rect 811 47 867 123
rect 897 89 953 177
rect 897 55 908 89
rect 942 55 953 89
rect 897 47 953 55
rect 983 157 1039 177
rect 983 123 994 157
rect 1028 123 1039 157
rect 983 47 1039 123
rect 1069 89 1126 177
rect 1069 55 1080 89
rect 1114 55 1126 89
rect 1069 47 1126 55
<< pdiff >>
rect 32 485 85 497
rect 32 451 40 485
rect 74 451 85 485
rect 32 417 85 451
rect 32 383 40 417
rect 74 383 85 417
rect 32 297 85 383
rect 115 477 171 497
rect 115 443 126 477
rect 160 443 171 477
rect 115 297 171 443
rect 201 485 257 497
rect 201 451 212 485
rect 246 451 257 485
rect 201 297 257 451
rect 287 477 343 497
rect 287 443 298 477
rect 332 443 343 477
rect 287 297 343 443
rect 373 405 429 497
rect 373 371 384 405
rect 418 371 429 405
rect 373 297 429 371
rect 459 489 515 497
rect 459 455 470 489
rect 504 455 515 489
rect 459 297 515 455
rect 545 405 601 497
rect 545 371 556 405
rect 590 371 601 405
rect 545 297 601 371
rect 631 489 687 497
rect 631 455 642 489
rect 676 455 687 489
rect 631 297 687 455
rect 717 489 781 497
rect 717 455 732 489
rect 766 455 781 489
rect 717 297 781 455
rect 811 477 867 497
rect 811 443 822 477
rect 856 443 867 477
rect 811 382 867 443
rect 811 348 822 382
rect 856 348 867 382
rect 811 297 867 348
rect 897 485 953 497
rect 897 451 908 485
rect 942 451 953 485
rect 897 297 953 451
rect 983 477 1039 497
rect 983 443 994 477
rect 1028 443 1039 477
rect 983 382 1039 443
rect 983 348 994 382
rect 1028 348 1039 382
rect 983 297 1039 348
rect 1069 485 1122 497
rect 1069 451 1080 485
rect 1114 451 1122 485
rect 1069 410 1122 451
rect 1069 376 1080 410
rect 1114 376 1122 410
rect 1069 297 1122 376
<< ndiffc >>
rect 40 123 74 157
rect 126 55 160 89
rect 212 123 246 157
rect 298 55 332 89
rect 384 123 418 157
rect 470 55 504 89
rect 556 123 590 157
rect 642 55 676 89
rect 736 91 770 125
rect 822 123 856 157
rect 908 55 942 89
rect 994 123 1028 157
rect 1080 55 1114 89
<< pdiffc >>
rect 40 451 74 485
rect 40 383 74 417
rect 126 443 160 477
rect 212 451 246 485
rect 298 443 332 477
rect 384 371 418 405
rect 470 455 504 489
rect 556 371 590 405
rect 642 455 676 489
rect 732 455 766 489
rect 822 443 856 477
rect 822 348 856 382
rect 908 451 942 485
rect 994 443 1028 477
rect 994 348 1028 382
rect 1080 451 1114 485
rect 1080 376 1114 410
<< poly >>
rect 85 497 115 523
rect 171 497 201 523
rect 257 497 287 523
rect 343 497 373 523
rect 429 497 459 523
rect 515 497 545 523
rect 601 497 631 523
rect 687 497 717 523
rect 781 497 811 523
rect 867 497 897 523
rect 953 497 983 523
rect 1039 497 1069 523
rect 85 265 115 297
rect 171 265 201 297
rect 257 265 287 297
rect 343 265 373 297
rect 429 265 459 297
rect 515 265 545 297
rect 601 265 631 297
rect 687 265 717 297
rect 781 265 811 297
rect 867 265 897 297
rect 953 265 983 297
rect 1039 265 1069 297
rect 25 249 295 265
rect 25 215 41 249
rect 75 215 109 249
rect 143 215 177 249
rect 211 215 245 249
rect 279 215 295 249
rect 25 199 295 215
rect 343 249 631 265
rect 343 215 415 249
rect 449 215 501 249
rect 535 215 581 249
rect 615 215 631 249
rect 343 199 631 215
rect 673 249 739 265
rect 673 215 689 249
rect 723 215 739 249
rect 673 199 739 215
rect 781 249 1069 265
rect 781 215 797 249
rect 831 215 865 249
rect 899 215 933 249
rect 967 215 1001 249
rect 1035 215 1069 249
rect 781 199 1069 215
rect 85 177 115 199
rect 171 177 201 199
rect 257 177 287 199
rect 343 177 373 199
rect 429 177 459 199
rect 515 177 545 199
rect 601 177 631 199
rect 695 177 725 199
rect 781 177 811 199
rect 867 177 897 199
rect 953 177 983 199
rect 1039 177 1069 199
rect 85 21 115 47
rect 171 21 201 47
rect 257 21 287 47
rect 343 21 373 47
rect 429 21 459 47
rect 515 21 545 47
rect 601 21 631 47
rect 695 21 725 47
rect 781 21 811 47
rect 867 21 897 47
rect 953 21 983 47
rect 1039 21 1069 47
<< polycont >>
rect 41 215 75 249
rect 109 215 143 249
rect 177 215 211 249
rect 245 215 279 249
rect 415 215 449 249
rect 501 215 535 249
rect 581 215 615 249
rect 689 215 723 249
rect 797 215 831 249
rect 865 215 899 249
rect 933 215 967 249
rect 1001 215 1035 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 24 485 81 527
rect 24 451 40 485
rect 74 451 81 485
rect 24 417 81 451
rect 24 383 40 417
rect 74 383 81 417
rect 115 477 162 493
rect 115 443 126 477
rect 160 443 162 477
rect 196 485 262 527
rect 196 451 212 485
rect 246 451 262 485
rect 296 489 692 493
rect 296 477 470 489
rect 115 417 162 443
rect 296 443 298 477
rect 332 455 470 477
rect 504 455 642 489
rect 676 455 692 489
rect 726 489 782 527
rect 726 455 732 489
rect 766 455 782 489
rect 332 443 334 455
rect 296 417 334 443
rect 726 439 782 455
rect 816 477 858 493
rect 816 443 822 477
rect 856 443 858 477
rect 892 485 958 527
rect 892 451 908 485
rect 942 451 958 485
rect 992 477 1030 493
rect 115 383 334 417
rect 816 417 858 443
rect 992 443 994 477
rect 1028 443 1030 477
rect 992 417 1030 443
rect 816 405 1030 417
rect 24 364 81 383
rect 368 371 384 405
rect 418 371 556 405
rect 590 382 1030 405
rect 590 371 822 382
rect 787 348 822 371
rect 856 348 994 382
rect 1028 348 1030 382
rect 1064 485 1130 527
rect 1064 451 1080 485
rect 1114 451 1130 485
rect 1064 410 1130 451
rect 1064 376 1080 410
rect 1114 376 1130 410
rect 787 340 1030 348
rect 115 303 739 337
rect 115 264 295 303
rect 25 249 295 264
rect 25 215 41 249
rect 75 215 109 249
rect 143 215 177 249
rect 211 215 245 249
rect 279 215 295 249
rect 25 203 295 215
rect 397 249 655 269
rect 397 215 415 249
rect 449 215 501 249
rect 535 215 581 249
rect 615 215 655 249
rect 397 214 655 215
rect 689 249 739 303
rect 787 289 1167 340
rect 723 215 739 249
rect 689 198 739 215
rect 781 249 1051 255
rect 781 215 797 249
rect 831 215 865 249
rect 899 215 933 249
rect 967 215 1001 249
rect 1035 215 1051 249
rect 781 203 1051 215
rect 1085 169 1167 289
rect 24 157 772 164
rect 24 123 40 157
rect 74 123 212 157
rect 246 123 384 157
rect 418 123 556 157
rect 590 125 772 157
rect 590 123 736 125
rect 726 91 736 123
rect 770 91 772 125
rect 806 157 1167 169
rect 806 123 822 157
rect 856 123 994 157
rect 1028 123 1167 157
rect 726 89 772 91
rect 110 55 126 89
rect 160 55 176 89
rect 110 17 176 55
rect 282 55 298 89
rect 332 55 348 89
rect 282 17 348 55
rect 454 55 470 89
rect 504 55 520 89
rect 454 17 520 55
rect 626 55 642 89
rect 676 55 692 89
rect 626 17 692 55
rect 726 55 908 89
rect 942 55 1080 89
rect 1114 55 1130 89
rect 726 51 1130 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
flabel locali s 1133 153 1167 187 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 857 221 891 255 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 397 221 431 255 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 213 289 247 323 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
rlabel comment s 0 0 0 0 4 o21ai_4
rlabel metal1 s 0 -48 1196 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1196 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1196 544
string GDS_END 1261856
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1253802
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 5.980 0.000 
<< end >>
