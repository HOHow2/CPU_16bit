magic
tech sky130A
magscale 1 2
timestamp 1738263620
<< nwell >>
rect -38 261 1970 582
<< pwell >>
rect 704 157 886 201
rect 1194 157 1931 203
rect 1 21 1931 157
rect 29 -17 63 21
<< locali >>
rect 18 195 88 325
rect 274 143 330 333
rect 1378 315 1444 484
rect 1378 299 1460 315
rect 1413 289 1460 299
rect 1422 173 1460 289
rect 1411 165 1460 173
rect 1380 148 1460 165
rect 1762 299 1829 493
rect 1380 61 1446 148
rect 1786 177 1829 299
rect 1778 53 1829 177
<< obsli1 >>
rect 0 527 1932 561
rect 35 393 69 493
rect 103 427 169 527
rect 35 359 168 393
rect 122 161 168 359
rect 35 127 168 161
rect 35 69 69 127
rect 103 17 169 93
rect 203 69 240 493
rect 288 435 341 527
rect 375 408 425 493
rect 467 438 688 472
rect 364 382 425 408
rect 364 161 398 382
rect 432 225 480 344
rect 514 331 620 404
rect 514 191 548 331
rect 654 315 688 438
rect 722 367 756 527
rect 790 427 840 493
rect 885 433 1062 467
rect 654 297 756 315
rect 364 135 409 161
rect 443 147 548 191
rect 582 263 756 297
rect 291 17 341 109
rect 375 107 409 135
rect 582 107 616 263
rect 722 249 756 263
rect 658 213 698 219
rect 790 213 824 427
rect 858 249 896 393
rect 658 153 824 213
rect 930 207 994 399
rect 375 73 442 107
rect 481 73 616 107
rect 680 17 754 117
rect 790 107 824 153
rect 901 141 994 207
rect 1028 265 1062 433
rect 1098 427 1161 527
rect 1208 381 1276 493
rect 1096 306 1276 381
rect 1310 325 1344 527
rect 1238 265 1276 306
rect 1478 344 1513 527
rect 1581 343 1647 489
rect 1028 199 1204 265
rect 1238 199 1388 265
rect 1028 107 1062 199
rect 1238 165 1278 199
rect 790 73 871 107
rect 905 73 1062 107
rect 1117 17 1159 123
rect 1212 60 1278 165
rect 1593 265 1647 343
rect 1685 299 1728 527
rect 1863 299 1913 527
rect 1593 199 1752 265
rect 1312 17 1346 139
rect 1593 123 1633 199
rect 1480 17 1514 120
rect 1581 69 1633 123
rect 1678 17 1744 165
rect 1863 17 1913 181
rect 0 -17 1932 17
<< metal1 >>
rect 0 496 1932 592
rect 0 -48 1932 48
<< obsm1 >>
rect 114 388 172 397
rect 534 388 592 397
rect 848 388 906 397
rect 114 360 906 388
rect 114 351 172 360
rect 534 351 592 360
rect 848 351 906 360
rect 193 320 251 329
rect 431 320 489 329
rect 935 320 993 329
rect 193 292 993 320
rect 193 283 251 292
rect 431 283 489 292
rect 935 283 993 292
<< labels >>
rlabel locali s 18 195 88 325 6 CLK
port 1 nsew clock input
rlabel locali s 274 143 330 333 6 D
port 2 nsew signal input
rlabel metal1 s 0 -48 1932 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1 21 1931 157 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1194 157 1931 203 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 704 157 886 201 6 VNB
port 4 nsew ground bidirectional
rlabel nwell s -38 261 1970 582 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 496 1932 592 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 1380 61 1446 148 6 Q
port 7 nsew signal output
rlabel locali s 1380 148 1460 165 6 Q
port 7 nsew signal output
rlabel locali s 1411 165 1460 173 6 Q
port 7 nsew signal output
rlabel locali s 1422 173 1460 289 6 Q
port 7 nsew signal output
rlabel locali s 1413 289 1460 299 6 Q
port 7 nsew signal output
rlabel locali s 1378 299 1460 315 6 Q
port 7 nsew signal output
rlabel locali s 1378 315 1444 484 6 Q
port 7 nsew signal output
rlabel locali s 1778 53 1829 177 6 Q_N
port 8 nsew signal output
rlabel locali s 1786 177 1829 299 6 Q_N
port 8 nsew signal output
rlabel locali s 1762 299 1829 493 6 Q_N
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1932 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2744370
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2729288
<< end >>
