magic
tech sky130A
magscale 1 2
timestamp 1738263620
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 458 163 735 203
rect 1 27 735 163
rect 29 -17 63 27
rect 461 21 735 27
<< scnmos >>
rect 79 53 109 137
rect 271 53 301 137
rect 343 53 373 137
rect 424 53 454 137
rect 543 47 573 177
rect 627 47 657 177
<< scpmoshvt >>
rect 79 311 109 395
rect 267 311 297 395
rect 351 311 381 395
rect 446 297 476 381
rect 543 297 573 497
rect 627 297 657 497
<< ndiff >>
rect 484 137 543 177
rect 27 99 79 137
rect 27 65 35 99
rect 69 65 79 99
rect 27 53 79 65
rect 109 111 165 137
rect 109 77 123 111
rect 157 77 165 111
rect 109 53 165 77
rect 219 111 271 137
rect 219 77 227 111
rect 261 77 271 111
rect 219 53 271 77
rect 301 53 343 137
rect 373 53 424 137
rect 454 116 543 137
rect 454 82 498 116
rect 532 82 543 116
rect 454 53 543 82
rect 487 47 543 53
rect 573 123 627 177
rect 573 89 583 123
rect 617 89 627 123
rect 573 47 627 89
rect 657 120 709 177
rect 657 86 667 120
rect 701 86 709 120
rect 657 47 709 86
<< pdiff >>
rect 491 477 543 497
rect 491 443 499 477
rect 533 443 543 477
rect 491 408 543 443
rect 27 365 79 395
rect 27 331 35 365
rect 69 331 79 365
rect 27 311 79 331
rect 109 365 161 395
rect 109 331 119 365
rect 153 331 161 365
rect 109 311 161 331
rect 215 369 267 395
rect 215 335 223 369
rect 257 335 267 369
rect 215 311 267 335
rect 297 387 351 395
rect 297 353 307 387
rect 341 353 351 387
rect 297 311 351 353
rect 381 381 431 395
rect 491 381 499 408
rect 381 362 446 381
rect 381 328 402 362
rect 436 328 446 362
rect 381 311 446 328
rect 396 297 446 311
rect 476 374 499 381
rect 533 374 543 408
rect 476 297 543 374
rect 573 477 627 497
rect 573 443 583 477
rect 617 443 627 477
rect 573 409 627 443
rect 573 375 583 409
rect 617 375 627 409
rect 573 297 627 375
rect 657 477 709 497
rect 657 443 667 477
rect 701 443 709 477
rect 657 409 709 443
rect 657 375 667 409
rect 701 375 709 409
rect 657 297 709 375
<< ndiffc >>
rect 35 65 69 99
rect 123 77 157 111
rect 227 77 261 111
rect 498 82 532 116
rect 583 89 617 123
rect 667 86 701 120
<< pdiffc >>
rect 499 443 533 477
rect 35 331 69 365
rect 119 331 153 365
rect 223 335 257 369
rect 307 353 341 387
rect 402 328 436 362
rect 499 374 533 408
rect 583 443 617 477
rect 583 375 617 409
rect 667 443 701 477
rect 667 375 701 409
<< poly >>
rect 351 477 407 500
rect 543 497 573 523
rect 627 497 657 523
rect 351 443 363 477
rect 397 443 407 477
rect 351 427 407 443
rect 79 395 109 425
rect 267 395 297 425
rect 351 395 381 427
rect 446 381 476 407
rect 79 265 109 311
rect 267 265 297 311
rect 28 259 109 265
rect 21 249 109 259
rect 21 215 37 249
rect 71 215 109 249
rect 21 205 109 215
rect 28 199 109 205
rect 217 249 301 265
rect 217 215 227 249
rect 261 215 301 249
rect 351 240 381 311
rect 446 265 476 297
rect 543 265 573 297
rect 627 265 657 297
rect 217 199 301 215
rect 79 137 109 199
rect 271 137 301 199
rect 343 203 381 240
rect 424 249 478 265
rect 424 215 434 249
rect 468 215 478 249
rect 343 137 373 203
rect 424 199 478 215
rect 520 249 657 265
rect 520 215 530 249
rect 564 215 657 249
rect 520 199 657 215
rect 424 137 454 199
rect 543 177 573 199
rect 627 177 657 199
rect 79 27 109 53
rect 271 27 301 53
rect 343 27 373 53
rect 424 27 454 53
rect 543 21 573 47
rect 627 21 657 47
<< polycont >>
rect 363 443 397 477
rect 37 215 71 249
rect 227 215 261 249
rect 434 215 468 249
rect 530 215 564 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 17 365 80 527
rect 206 426 329 527
rect 17 331 35 365
rect 69 331 80 365
rect 17 315 80 331
rect 116 365 171 381
rect 116 331 119 365
rect 153 331 171 365
rect 29 249 82 265
rect 29 215 37 249
rect 71 215 82 249
rect 29 149 82 215
rect 116 249 171 331
rect 210 369 257 392
rect 210 335 223 369
rect 291 391 329 426
rect 363 477 458 493
rect 397 443 458 477
rect 363 425 458 443
rect 492 477 535 527
rect 492 443 499 477
rect 533 443 535 477
rect 492 408 535 443
rect 291 387 357 391
rect 291 353 307 387
rect 341 353 357 387
rect 402 362 440 378
rect 210 319 257 335
rect 436 328 440 362
rect 492 374 499 408
rect 533 374 535 408
rect 492 358 535 374
rect 575 477 632 493
rect 575 443 583 477
rect 617 443 632 477
rect 575 409 632 443
rect 575 375 583 409
rect 617 375 632 409
rect 575 359 632 375
rect 402 319 440 328
rect 210 285 564 319
rect 116 215 227 249
rect 261 215 283 249
rect 116 203 283 215
rect 17 99 71 115
rect 17 65 35 99
rect 69 65 71 99
rect 17 17 71 65
rect 116 111 171 203
rect 317 114 368 285
rect 518 249 564 285
rect 116 77 123 111
rect 157 77 171 111
rect 116 61 171 77
rect 211 111 368 114
rect 211 77 227 111
rect 261 77 368 111
rect 211 61 368 77
rect 402 215 434 249
rect 468 215 484 249
rect 402 153 484 215
rect 518 215 530 249
rect 518 199 564 215
rect 598 289 632 359
rect 666 477 719 527
rect 666 443 667 477
rect 701 443 719 477
rect 666 409 719 443
rect 666 375 667 409
rect 701 375 719 409
rect 666 325 719 375
rect 598 185 719 289
rect 402 61 444 153
rect 598 143 632 185
rect 583 123 632 143
rect 482 82 498 116
rect 532 82 548 116
rect 482 17 548 82
rect 617 89 632 123
rect 583 51 632 89
rect 666 120 719 149
rect 666 86 667 120
rect 701 86 719 120
rect 666 17 719 86
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel locali s 402 425 436 459 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel locali s 584 85 618 119 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 584 425 618 459 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 29 221 63 255 0 FreeSans 400 0 0 0 A_N
port 1 nsew signal input
flabel locali s 402 153 436 187 0 FreeSans 400 0 0 0 C
port 3 nsew signal input
flabel locali s 672 221 706 255 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 and3b_2
rlabel metal1 s 0 -48 736 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 736 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_END 3082846
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3076298
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
