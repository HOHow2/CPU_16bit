magic
tech sky130A
magscale 1 2
timestamp 1738263620
<< nwell >>
rect -38 261 2062 582
<< pwell >>
rect 1 21 2023 203
rect 30 -17 64 21
<< locali >>
rect 22 261 66 393
rect 103 349 169 417
rect 271 349 337 417
rect 395 349 505 417
rect 607 349 673 417
rect 103 315 673 349
rect 22 215 350 261
rect 395 198 473 315
rect 517 199 711 265
rect 755 215 1093 257
rect 1219 215 1539 260
rect 1659 215 1997 256
rect 439 161 473 198
rect 439 127 1113 161
rect 1961 151 1997 215
<< obsli1 >>
rect 0 527 2024 561
rect 19 451 741 485
rect 707 349 741 451
rect 779 383 845 527
rect 879 349 913 493
rect 954 383 1088 527
rect 1128 349 1162 493
rect 1243 383 1309 527
rect 1343 349 1377 493
rect 1411 383 1477 527
rect 1511 349 1545 493
rect 1683 383 1749 527
rect 1783 349 1817 493
rect 1851 383 1917 527
rect 1951 349 1985 493
rect 707 315 1985 349
rect 35 127 405 161
rect 1243 127 1901 161
rect 35 51 69 127
rect 103 17 169 93
rect 203 51 237 127
rect 371 93 405 127
rect 271 17 337 93
rect 371 59 757 93
rect 795 59 1561 93
rect 1599 17 1665 93
rect 1699 51 1733 127
rect 1767 17 1833 93
rect 1867 51 1901 127
rect 1937 17 2005 93
rect 0 -17 2024 17
<< metal1 >>
rect 0 496 2024 592
rect 0 -48 2024 48
<< labels >>
rlabel locali s 755 215 1093 257 6 A1
port 1 nsew signal input
rlabel locali s 1219 215 1539 260 6 A2
port 2 nsew signal input
rlabel locali s 1961 151 1997 215 6 A3
port 3 nsew signal input
rlabel locali s 1659 215 1997 256 6 A3
port 3 nsew signal input
rlabel locali s 517 199 711 265 6 B1
port 4 nsew signal input
rlabel locali s 22 215 350 261 6 B2
port 5 nsew signal input
rlabel locali s 22 261 66 393 6 B2
port 5 nsew signal input
rlabel metal1 s 0 -48 2024 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 1 21 2023 203 6 VNB
port 7 nsew ground bidirectional
rlabel nwell s -38 261 2062 582 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 496 2024 592 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 439 127 1113 161 6 Y
port 10 nsew signal output
rlabel locali s 439 161 473 198 6 Y
port 10 nsew signal output
rlabel locali s 395 198 473 315 6 Y
port 10 nsew signal output
rlabel locali s 103 315 673 349 6 Y
port 10 nsew signal output
rlabel locali s 607 349 673 417 6 Y
port 10 nsew signal output
rlabel locali s 395 349 505 417 6 Y
port 10 nsew signal output
rlabel locali s 271 349 337 417 6 Y
port 10 nsew signal output
rlabel locali s 103 349 169 417 6 Y
port 10 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2024 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3578196
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3562022
<< end >>
