magic
tech sky130A
magscale 1 2
timestamp 1738263620
<< nwell >>
rect -38 261 498 582
<< pwell >>
rect 98 157 459 203
rect 1 21 459 157
rect 30 -17 64 21
<< locali >>
rect 324 425 443 493
rect 17 199 109 345
rect 324 161 359 425
rect 395 195 443 391
rect 324 51 443 161
<< obsli1 >>
rect 0 527 460 561
rect 17 413 69 493
rect 103 447 290 527
rect 17 379 290 413
rect 143 165 290 379
rect 17 131 290 165
rect 17 51 69 131
rect 103 17 290 97
rect 0 -17 460 17
<< metal1 >>
rect 0 496 460 592
rect 0 -48 460 48
<< labels >>
rlabel locali s 395 195 443 391 6 A
port 1 nsew signal input
rlabel locali s 17 199 109 345 6 TE
port 2 nsew signal input
rlabel metal1 s 0 -48 460 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1 21 459 157 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 98 157 459 203 6 VNB
port 4 nsew ground bidirectional
rlabel nwell s -38 261 498 582 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 496 460 592 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 324 51 443 161 6 Z
port 7 nsew signal output
rlabel locali s 324 161 359 425 6 Z
port 7 nsew signal output
rlabel locali s 324 425 443 493 6 Z
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 460 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2096840
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2092328
<< end >>
